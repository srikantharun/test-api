// (C) Copyright 2024 Axelera AI B.V.
// All Rights Reserved
// *** Axelera AI Confidential ***
//
// Description: NOC Top
// Owners: Joao Martins <joao.martins@axelera.ai>
//         Deeptanshu Sekhri <deeptanshu.sekhri@axelera.ai>
//         Tasos Psarras <anastasios.psarras@axelera.ai>


module noc_top (
    input wire                              i_ref_clk,
    // DFT Interface
    input  logic                            test_mode,
    input  logic                            scan_en,
    // SDMA0
    input wire                              i_sdma_0_clk,
    input wire                              i_sdma_0_ao_rst_n,
    input wire                              i_sdma_0_global_rst_n,
    output logic[sdma_pkg::NUM_CHNLS-1:0]   o_sdma_0_int,
    input logic                             i_sdma_0_clock_throttle,
    // SDMA1
    input wire                              i_sdma_1_clk,
    input wire                              i_sdma_1_ao_rst_n,
    input wire                              i_sdma_1_global_rst_n,
    output logic[sdma_pkg::NUM_CHNLS-1:0]   o_sdma_1_int,
    input logic                             i_sdma_1_clock_throttle,
    input  logic                            i_sdma_inter_core_sync,
    // rest
    output logic[15:0]                                         o_obs,
    output logic                                               o_irq,
    input  wire                                                i_aic_0_aon_clk,
    input  wire                                                i_aic_0_aon_rst_n,
    input  wire                                                i_aic_0_clk,
    input  wire                                                i_aic_0_clken,
    input  chip_pkg::chip_axi_addr_t                           i_aic_0_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_0_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_0_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_0_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_0_init_ht_axi_s_arlen,
    input  logic                                               i_aic_0_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_0_init_ht_axi_s_arprot,
    output logic                                               o_aic_0_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_0_init_ht_axi_s_arsize,
    input  logic                                               i_aic_0_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_aic_0_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_0_init_ht_axi_s_rid,
    output logic                                               o_aic_0_init_ht_axi_s_rlast,
    input  logic                                               i_aic_0_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_0_init_ht_axi_s_rresp,
    output logic                                               o_aic_0_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_0_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_0_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_0_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_0_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_0_init_ht_axi_s_awlen,
    input  logic                                               i_aic_0_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_0_init_ht_axi_s_awprot,
    output logic                                               o_aic_0_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_0_init_ht_axi_s_awsize,
    input  logic                                               i_aic_0_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_0_init_ht_axi_s_bid,
    input  logic                                               i_aic_0_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_0_init_ht_axi_s_bresp,
    output logic                                               o_aic_0_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_aic_0_init_ht_axi_s_wdata,
    input  logic                                               i_aic_0_init_ht_axi_s_wlast,
    output logic                                               o_aic_0_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_aic_0_init_ht_axi_s_wstrb,
    input  logic                                               i_aic_0_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_0_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_0_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_0_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_0_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_0_init_lt_axi_s_arlen,
    input  logic                                               i_aic_0_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_0_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_aic_0_init_lt_axi_s_arqos,
    output logic                                               o_aic_0_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_0_init_lt_axi_s_arsize,
    input  logic                                               i_aic_0_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_0_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_0_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_0_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_0_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_0_init_lt_axi_s_awlen,
    input  logic                                               i_aic_0_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_0_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_aic_0_init_lt_axi_s_awqos,
    output logic                                               o_aic_0_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_0_init_lt_axi_s_awsize,
    input  logic                                               i_aic_0_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_0_init_lt_axi_s_bid,
    input  logic                                               i_aic_0_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_0_init_lt_axi_s_bresp,
    output logic                                               o_aic_0_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_0_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_0_init_lt_axi_s_rid,
    output logic                                               o_aic_0_init_lt_axi_s_rlast,
    input  logic                                               i_aic_0_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_0_init_lt_axi_s_rresp,
    output logic                                               o_aic_0_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_0_init_lt_axi_s_wdata,
    input  logic                                               i_aic_0_init_lt_axi_s_wlast,
    output logic                                               o_aic_0_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_aic_0_init_lt_axi_s_wstrb,
    input  logic                                               i_aic_0_init_lt_axi_s_wvalid,
    output logic                                               o_aic_0_pwr_idle_val,
    output logic                                               o_aic_0_pwr_idle_ack,
    input  logic                                               i_aic_0_pwr_idle_req,
    input  wire                                                i_aic_0_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_aic_0_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_aic_0_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_aic_0_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_0_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_aic_0_targ_lt_axi_m_arlen,
    output logic                                               o_aic_0_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_aic_0_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_aic_0_targ_lt_axi_m_arqos,
    input  logic                                               i_aic_0_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_aic_0_targ_lt_axi_m_arsize,
    output logic                                               o_aic_0_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_aic_0_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_aic_0_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_aic_0_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_0_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_aic_0_targ_lt_axi_m_awlen,
    output logic                                               o_aic_0_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_aic_0_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_aic_0_targ_lt_axi_m_awqos,
    input  logic                                               i_aic_0_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_aic_0_targ_lt_axi_m_awsize,
    output logic                                               o_aic_0_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_0_targ_lt_axi_m_bid,
    output logic                                               o_aic_0_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_aic_0_targ_lt_axi_m_bresp,
    input  logic                                               i_aic_0_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_0_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_0_targ_lt_axi_m_rid,
    input  logic                                               i_aic_0_targ_lt_axi_m_rlast,
    output logic                                               o_aic_0_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_aic_0_targ_lt_axi_m_rresp,
    input  logic                                               i_aic_0_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_0_targ_lt_axi_m_wdata,
    output logic                                               o_aic_0_targ_lt_axi_m_wlast,
    input  logic                                               i_aic_0_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_aic_0_targ_lt_axi_m_wstrb,
    output logic                                               o_aic_0_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_aic_0_targ_syscfg_apb_m_paddr,
    output logic                                               o_aic_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_aic_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_aic_0_targ_syscfg_apb_m_prdata,
    input  logic                                               i_aic_0_targ_syscfg_apb_m_pready,
    output logic                                               o_aic_0_targ_syscfg_apb_m_psel,
    input  logic                                               i_aic_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_aic_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_aic_0_targ_syscfg_apb_m_pwdata,
    output logic                                               o_aic_0_targ_syscfg_apb_m_pwrite,
    output logic                                               o_aic_0_pwr_tok_idle_val,
    output logic                                               o_aic_0_pwr_tok_idle_ack,
    input  logic                                               i_aic_0_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_aic_0_init_tok_ocpl_s_maddr,
    input  logic                                               i_aic_0_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_aic_0_init_tok_ocpl_s_mdata,
    output logic                                               o_aic_0_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_aic_0_targ_tok_ocpl_m_maddr,
    output logic                                               o_aic_0_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_aic_0_targ_tok_ocpl_m_mdata,
    input  logic                                               i_aic_0_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_aic_1_aon_clk,
    input  wire                                                i_aic_1_aon_rst_n,
    input  wire                                                i_aic_1_clk,
    input  wire                                                i_aic_1_clken,
    input  chip_pkg::chip_axi_addr_t                           i_aic_1_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_1_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_1_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_1_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_1_init_ht_axi_s_arlen,
    input  logic                                               i_aic_1_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_1_init_ht_axi_s_arprot,
    output logic                                               o_aic_1_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_1_init_ht_axi_s_arsize,
    input  logic                                               i_aic_1_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_aic_1_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_1_init_ht_axi_s_rid,
    output logic                                               o_aic_1_init_ht_axi_s_rlast,
    input  logic                                               i_aic_1_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_1_init_ht_axi_s_rresp,
    output logic                                               o_aic_1_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_1_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_1_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_1_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_1_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_1_init_ht_axi_s_awlen,
    input  logic                                               i_aic_1_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_1_init_ht_axi_s_awprot,
    output logic                                               o_aic_1_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_1_init_ht_axi_s_awsize,
    input  logic                                               i_aic_1_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_1_init_ht_axi_s_bid,
    input  logic                                               i_aic_1_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_1_init_ht_axi_s_bresp,
    output logic                                               o_aic_1_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_aic_1_init_ht_axi_s_wdata,
    input  logic                                               i_aic_1_init_ht_axi_s_wlast,
    output logic                                               o_aic_1_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_aic_1_init_ht_axi_s_wstrb,
    input  logic                                               i_aic_1_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_1_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_1_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_1_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_1_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_1_init_lt_axi_s_arlen,
    input  logic                                               i_aic_1_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_1_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_aic_1_init_lt_axi_s_arqos,
    output logic                                               o_aic_1_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_1_init_lt_axi_s_arsize,
    input  logic                                               i_aic_1_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_1_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_1_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_1_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_1_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_1_init_lt_axi_s_awlen,
    input  logic                                               i_aic_1_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_1_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_aic_1_init_lt_axi_s_awqos,
    output logic                                               o_aic_1_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_1_init_lt_axi_s_awsize,
    input  logic                                               i_aic_1_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_1_init_lt_axi_s_bid,
    input  logic                                               i_aic_1_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_1_init_lt_axi_s_bresp,
    output logic                                               o_aic_1_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_1_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_1_init_lt_axi_s_rid,
    output logic                                               o_aic_1_init_lt_axi_s_rlast,
    input  logic                                               i_aic_1_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_1_init_lt_axi_s_rresp,
    output logic                                               o_aic_1_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_1_init_lt_axi_s_wdata,
    input  logic                                               i_aic_1_init_lt_axi_s_wlast,
    output logic                                               o_aic_1_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_aic_1_init_lt_axi_s_wstrb,
    input  logic                                               i_aic_1_init_lt_axi_s_wvalid,
    output logic                                               o_aic_1_pwr_idle_val,
    output logic                                               o_aic_1_pwr_idle_ack,
    input  logic                                               i_aic_1_pwr_idle_req,
    input  wire                                                i_aic_1_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_aic_1_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_aic_1_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_aic_1_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_1_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_aic_1_targ_lt_axi_m_arlen,
    output logic                                               o_aic_1_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_aic_1_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_aic_1_targ_lt_axi_m_arqos,
    input  logic                                               i_aic_1_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_aic_1_targ_lt_axi_m_arsize,
    output logic                                               o_aic_1_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_aic_1_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_aic_1_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_aic_1_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_1_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_aic_1_targ_lt_axi_m_awlen,
    output logic                                               o_aic_1_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_aic_1_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_aic_1_targ_lt_axi_m_awqos,
    input  logic                                               i_aic_1_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_aic_1_targ_lt_axi_m_awsize,
    output logic                                               o_aic_1_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_1_targ_lt_axi_m_bid,
    output logic                                               o_aic_1_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_aic_1_targ_lt_axi_m_bresp,
    input  logic                                               i_aic_1_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_1_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_1_targ_lt_axi_m_rid,
    input  logic                                               i_aic_1_targ_lt_axi_m_rlast,
    output logic                                               o_aic_1_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_aic_1_targ_lt_axi_m_rresp,
    input  logic                                               i_aic_1_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_1_targ_lt_axi_m_wdata,
    output logic                                               o_aic_1_targ_lt_axi_m_wlast,
    input  logic                                               i_aic_1_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_aic_1_targ_lt_axi_m_wstrb,
    output logic                                               o_aic_1_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_aic_1_targ_syscfg_apb_m_paddr,
    output logic                                               o_aic_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_aic_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_aic_1_targ_syscfg_apb_m_prdata,
    input  logic                                               i_aic_1_targ_syscfg_apb_m_pready,
    output logic                                               o_aic_1_targ_syscfg_apb_m_psel,
    input  logic                                               i_aic_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_aic_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_aic_1_targ_syscfg_apb_m_pwdata,
    output logic                                               o_aic_1_targ_syscfg_apb_m_pwrite,
    output logic                                               o_aic_1_pwr_tok_idle_val,
    output logic                                               o_aic_1_pwr_tok_idle_ack,
    input  logic                                               i_aic_1_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_aic_1_init_tok_ocpl_s_maddr,
    input  logic                                               i_aic_1_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_aic_1_init_tok_ocpl_s_mdata,
    output logic                                               o_aic_1_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_aic_1_targ_tok_ocpl_m_maddr,
    output logic                                               o_aic_1_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_aic_1_targ_tok_ocpl_m_mdata,
    input  logic                                               i_aic_1_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_aic_2_aon_clk,
    input  wire                                                i_aic_2_aon_rst_n,
    input  wire                                                i_aic_2_clk,
    input  wire                                                i_aic_2_clken,
    input  chip_pkg::chip_axi_addr_t                           i_aic_2_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_2_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_2_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_2_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_2_init_ht_axi_s_arlen,
    input  logic                                               i_aic_2_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_2_init_ht_axi_s_arprot,
    output logic                                               o_aic_2_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_2_init_ht_axi_s_arsize,
    input  logic                                               i_aic_2_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_aic_2_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_2_init_ht_axi_s_rid,
    output logic                                               o_aic_2_init_ht_axi_s_rlast,
    input  logic                                               i_aic_2_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_2_init_ht_axi_s_rresp,
    output logic                                               o_aic_2_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_2_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_2_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_2_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_2_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_2_init_ht_axi_s_awlen,
    input  logic                                               i_aic_2_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_2_init_ht_axi_s_awprot,
    output logic                                               o_aic_2_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_2_init_ht_axi_s_awsize,
    input  logic                                               i_aic_2_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_2_init_ht_axi_s_bid,
    input  logic                                               i_aic_2_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_2_init_ht_axi_s_bresp,
    output logic                                               o_aic_2_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_aic_2_init_ht_axi_s_wdata,
    input  logic                                               i_aic_2_init_ht_axi_s_wlast,
    output logic                                               o_aic_2_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_aic_2_init_ht_axi_s_wstrb,
    input  logic                                               i_aic_2_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_2_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_2_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_2_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_2_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_2_init_lt_axi_s_arlen,
    input  logic                                               i_aic_2_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_2_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_aic_2_init_lt_axi_s_arqos,
    output logic                                               o_aic_2_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_2_init_lt_axi_s_arsize,
    input  logic                                               i_aic_2_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_2_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_2_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_2_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_2_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_2_init_lt_axi_s_awlen,
    input  logic                                               i_aic_2_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_2_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_aic_2_init_lt_axi_s_awqos,
    output logic                                               o_aic_2_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_2_init_lt_axi_s_awsize,
    input  logic                                               i_aic_2_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_2_init_lt_axi_s_bid,
    input  logic                                               i_aic_2_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_2_init_lt_axi_s_bresp,
    output logic                                               o_aic_2_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_2_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_2_init_lt_axi_s_rid,
    output logic                                               o_aic_2_init_lt_axi_s_rlast,
    input  logic                                               i_aic_2_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_2_init_lt_axi_s_rresp,
    output logic                                               o_aic_2_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_2_init_lt_axi_s_wdata,
    input  logic                                               i_aic_2_init_lt_axi_s_wlast,
    output logic                                               o_aic_2_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_aic_2_init_lt_axi_s_wstrb,
    input  logic                                               i_aic_2_init_lt_axi_s_wvalid,
    output logic                                               o_aic_2_pwr_idle_val,
    output logic                                               o_aic_2_pwr_idle_ack,
    input  logic                                               i_aic_2_pwr_idle_req,
    input  wire                                                i_aic_2_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_aic_2_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_aic_2_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_aic_2_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_2_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_aic_2_targ_lt_axi_m_arlen,
    output logic                                               o_aic_2_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_aic_2_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_aic_2_targ_lt_axi_m_arqos,
    input  logic                                               i_aic_2_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_aic_2_targ_lt_axi_m_arsize,
    output logic                                               o_aic_2_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_aic_2_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_aic_2_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_aic_2_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_2_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_aic_2_targ_lt_axi_m_awlen,
    output logic                                               o_aic_2_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_aic_2_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_aic_2_targ_lt_axi_m_awqos,
    input  logic                                               i_aic_2_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_aic_2_targ_lt_axi_m_awsize,
    output logic                                               o_aic_2_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_2_targ_lt_axi_m_bid,
    output logic                                               o_aic_2_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_aic_2_targ_lt_axi_m_bresp,
    input  logic                                               i_aic_2_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_2_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_2_targ_lt_axi_m_rid,
    input  logic                                               i_aic_2_targ_lt_axi_m_rlast,
    output logic                                               o_aic_2_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_aic_2_targ_lt_axi_m_rresp,
    input  logic                                               i_aic_2_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_2_targ_lt_axi_m_wdata,
    output logic                                               o_aic_2_targ_lt_axi_m_wlast,
    input  logic                                               i_aic_2_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_aic_2_targ_lt_axi_m_wstrb,
    output logic                                               o_aic_2_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_aic_2_targ_syscfg_apb_m_paddr,
    output logic                                               o_aic_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_aic_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_aic_2_targ_syscfg_apb_m_prdata,
    input  logic                                               i_aic_2_targ_syscfg_apb_m_pready,
    output logic                                               o_aic_2_targ_syscfg_apb_m_psel,
    input  logic                                               i_aic_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_aic_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_aic_2_targ_syscfg_apb_m_pwdata,
    output logic                                               o_aic_2_targ_syscfg_apb_m_pwrite,
    output logic                                               o_aic_2_pwr_tok_idle_val,
    output logic                                               o_aic_2_pwr_tok_idle_ack,
    input  logic                                               i_aic_2_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_aic_2_init_tok_ocpl_s_maddr,
    input  logic                                               i_aic_2_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_aic_2_init_tok_ocpl_s_mdata,
    output logic                                               o_aic_2_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_aic_2_targ_tok_ocpl_m_maddr,
    output logic                                               o_aic_2_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_aic_2_targ_tok_ocpl_m_mdata,
    input  logic                                               i_aic_2_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_aic_3_aon_clk,
    input  wire                                                i_aic_3_aon_rst_n,
    input  wire                                                i_aic_3_clk,
    input  wire                                                i_aic_3_clken,
    input  chip_pkg::chip_axi_addr_t                           i_aic_3_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_3_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_3_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_3_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_3_init_ht_axi_s_arlen,
    input  logic                                               i_aic_3_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_3_init_ht_axi_s_arprot,
    output logic                                               o_aic_3_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_3_init_ht_axi_s_arsize,
    input  logic                                               i_aic_3_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_aic_3_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_3_init_ht_axi_s_rid,
    output logic                                               o_aic_3_init_ht_axi_s_rlast,
    input  logic                                               i_aic_3_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_3_init_ht_axi_s_rresp,
    output logic                                               o_aic_3_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_3_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_3_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_3_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_3_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_3_init_ht_axi_s_awlen,
    input  logic                                               i_aic_3_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_3_init_ht_axi_s_awprot,
    output logic                                               o_aic_3_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_3_init_ht_axi_s_awsize,
    input  logic                                               i_aic_3_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_3_init_ht_axi_s_bid,
    input  logic                                               i_aic_3_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_3_init_ht_axi_s_bresp,
    output logic                                               o_aic_3_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_aic_3_init_ht_axi_s_wdata,
    input  logic                                               i_aic_3_init_ht_axi_s_wlast,
    output logic                                               o_aic_3_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_aic_3_init_ht_axi_s_wstrb,
    input  logic                                               i_aic_3_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_3_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_3_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_3_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_3_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_3_init_lt_axi_s_arlen,
    input  logic                                               i_aic_3_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_3_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_aic_3_init_lt_axi_s_arqos,
    output logic                                               o_aic_3_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_3_init_lt_axi_s_arsize,
    input  logic                                               i_aic_3_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_3_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_3_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_3_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_3_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_3_init_lt_axi_s_awlen,
    input  logic                                               i_aic_3_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_3_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_aic_3_init_lt_axi_s_awqos,
    output logic                                               o_aic_3_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_3_init_lt_axi_s_awsize,
    input  logic                                               i_aic_3_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_3_init_lt_axi_s_bid,
    input  logic                                               i_aic_3_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_3_init_lt_axi_s_bresp,
    output logic                                               o_aic_3_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_3_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_3_init_lt_axi_s_rid,
    output logic                                               o_aic_3_init_lt_axi_s_rlast,
    input  logic                                               i_aic_3_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_3_init_lt_axi_s_rresp,
    output logic                                               o_aic_3_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_3_init_lt_axi_s_wdata,
    input  logic                                               i_aic_3_init_lt_axi_s_wlast,
    output logic                                               o_aic_3_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_aic_3_init_lt_axi_s_wstrb,
    input  logic                                               i_aic_3_init_lt_axi_s_wvalid,
    output logic                                               o_aic_3_pwr_idle_val,
    output logic                                               o_aic_3_pwr_idle_ack,
    input  logic                                               i_aic_3_pwr_idle_req,
    input  wire                                                i_aic_3_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_aic_3_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_aic_3_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_aic_3_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_3_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_aic_3_targ_lt_axi_m_arlen,
    output logic                                               o_aic_3_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_aic_3_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_aic_3_targ_lt_axi_m_arqos,
    input  logic                                               i_aic_3_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_aic_3_targ_lt_axi_m_arsize,
    output logic                                               o_aic_3_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_aic_3_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_aic_3_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_aic_3_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_3_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_aic_3_targ_lt_axi_m_awlen,
    output logic                                               o_aic_3_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_aic_3_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_aic_3_targ_lt_axi_m_awqos,
    input  logic                                               i_aic_3_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_aic_3_targ_lt_axi_m_awsize,
    output logic                                               o_aic_3_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_3_targ_lt_axi_m_bid,
    output logic                                               o_aic_3_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_aic_3_targ_lt_axi_m_bresp,
    input  logic                                               i_aic_3_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_3_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_3_targ_lt_axi_m_rid,
    input  logic                                               i_aic_3_targ_lt_axi_m_rlast,
    output logic                                               o_aic_3_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_aic_3_targ_lt_axi_m_rresp,
    input  logic                                               i_aic_3_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_3_targ_lt_axi_m_wdata,
    output logic                                               o_aic_3_targ_lt_axi_m_wlast,
    input  logic                                               i_aic_3_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_aic_3_targ_lt_axi_m_wstrb,
    output logic                                               o_aic_3_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_aic_3_targ_syscfg_apb_m_paddr,
    output logic                                               o_aic_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_aic_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_aic_3_targ_syscfg_apb_m_prdata,
    input  logic                                               i_aic_3_targ_syscfg_apb_m_pready,
    output logic                                               o_aic_3_targ_syscfg_apb_m_psel,
    input  logic                                               i_aic_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_aic_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_aic_3_targ_syscfg_apb_m_pwdata,
    output logic                                               o_aic_3_targ_syscfg_apb_m_pwrite,
    output logic                                               o_aic_3_pwr_tok_idle_val,
    output logic                                               o_aic_3_pwr_tok_idle_ack,
    input  logic                                               i_aic_3_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_aic_3_init_tok_ocpl_s_maddr,
    input  logic                                               i_aic_3_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_aic_3_init_tok_ocpl_s_mdata,
    output logic                                               o_aic_3_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_aic_3_targ_tok_ocpl_m_maddr,
    output logic                                               o_aic_3_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_aic_3_targ_tok_ocpl_m_mdata,
    input  logic                                               i_aic_3_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_aic_4_aon_clk,
    input  wire                                                i_aic_4_aon_rst_n,
    input  wire                                                i_aic_4_clk,
    input  wire                                                i_aic_4_clken,
    input  chip_pkg::chip_axi_addr_t                           i_aic_4_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_4_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_4_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_4_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_4_init_ht_axi_s_arlen,
    input  logic                                               i_aic_4_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_4_init_ht_axi_s_arprot,
    output logic                                               o_aic_4_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_4_init_ht_axi_s_arsize,
    input  logic                                               i_aic_4_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_aic_4_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_4_init_ht_axi_s_rid,
    output logic                                               o_aic_4_init_ht_axi_s_rlast,
    input  logic                                               i_aic_4_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_4_init_ht_axi_s_rresp,
    output logic                                               o_aic_4_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_4_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_4_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_4_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_4_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_4_init_ht_axi_s_awlen,
    input  logic                                               i_aic_4_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_4_init_ht_axi_s_awprot,
    output logic                                               o_aic_4_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_4_init_ht_axi_s_awsize,
    input  logic                                               i_aic_4_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_4_init_ht_axi_s_bid,
    input  logic                                               i_aic_4_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_4_init_ht_axi_s_bresp,
    output logic                                               o_aic_4_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_aic_4_init_ht_axi_s_wdata,
    input  logic                                               i_aic_4_init_ht_axi_s_wlast,
    output logic                                               o_aic_4_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_aic_4_init_ht_axi_s_wstrb,
    input  logic                                               i_aic_4_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_4_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_4_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_4_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_4_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_4_init_lt_axi_s_arlen,
    input  logic                                               i_aic_4_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_4_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_aic_4_init_lt_axi_s_arqos,
    output logic                                               o_aic_4_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_4_init_lt_axi_s_arsize,
    input  logic                                               i_aic_4_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_4_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_4_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_4_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_4_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_4_init_lt_axi_s_awlen,
    input  logic                                               i_aic_4_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_4_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_aic_4_init_lt_axi_s_awqos,
    output logic                                               o_aic_4_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_4_init_lt_axi_s_awsize,
    input  logic                                               i_aic_4_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_4_init_lt_axi_s_bid,
    input  logic                                               i_aic_4_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_4_init_lt_axi_s_bresp,
    output logic                                               o_aic_4_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_4_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_4_init_lt_axi_s_rid,
    output logic                                               o_aic_4_init_lt_axi_s_rlast,
    input  logic                                               i_aic_4_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_4_init_lt_axi_s_rresp,
    output logic                                               o_aic_4_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_4_init_lt_axi_s_wdata,
    input  logic                                               i_aic_4_init_lt_axi_s_wlast,
    output logic                                               o_aic_4_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_aic_4_init_lt_axi_s_wstrb,
    input  logic                                               i_aic_4_init_lt_axi_s_wvalid,
    output logic                                               o_aic_4_pwr_idle_val,
    output logic                                               o_aic_4_pwr_idle_ack,
    input  logic                                               i_aic_4_pwr_idle_req,
    input  wire                                                i_aic_4_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_aic_4_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_aic_4_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_aic_4_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_4_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_aic_4_targ_lt_axi_m_arlen,
    output logic                                               o_aic_4_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_aic_4_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_aic_4_targ_lt_axi_m_arqos,
    input  logic                                               i_aic_4_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_aic_4_targ_lt_axi_m_arsize,
    output logic                                               o_aic_4_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_aic_4_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_aic_4_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_aic_4_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_4_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_aic_4_targ_lt_axi_m_awlen,
    output logic                                               o_aic_4_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_aic_4_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_aic_4_targ_lt_axi_m_awqos,
    input  logic                                               i_aic_4_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_aic_4_targ_lt_axi_m_awsize,
    output logic                                               o_aic_4_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_4_targ_lt_axi_m_bid,
    output logic                                               o_aic_4_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_aic_4_targ_lt_axi_m_bresp,
    input  logic                                               i_aic_4_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_4_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_4_targ_lt_axi_m_rid,
    input  logic                                               i_aic_4_targ_lt_axi_m_rlast,
    output logic                                               o_aic_4_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_aic_4_targ_lt_axi_m_rresp,
    input  logic                                               i_aic_4_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_4_targ_lt_axi_m_wdata,
    output logic                                               o_aic_4_targ_lt_axi_m_wlast,
    input  logic                                               i_aic_4_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_aic_4_targ_lt_axi_m_wstrb,
    output logic                                               o_aic_4_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_aic_4_targ_syscfg_apb_m_paddr,
    output logic                                               o_aic_4_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_aic_4_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_aic_4_targ_syscfg_apb_m_prdata,
    input  logic                                               i_aic_4_targ_syscfg_apb_m_pready,
    output logic                                               o_aic_4_targ_syscfg_apb_m_psel,
    input  logic                                               i_aic_4_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_aic_4_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_aic_4_targ_syscfg_apb_m_pwdata,
    output logic                                               o_aic_4_targ_syscfg_apb_m_pwrite,
    output logic                                               o_aic_4_pwr_tok_idle_val,
    output logic                                               o_aic_4_pwr_tok_idle_ack,
    input  logic                                               i_aic_4_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_aic_4_init_tok_ocpl_s_maddr,
    input  logic                                               i_aic_4_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_aic_4_init_tok_ocpl_s_mdata,
    output logic                                               o_aic_4_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_aic_4_targ_tok_ocpl_m_maddr,
    output logic                                               o_aic_4_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_aic_4_targ_tok_ocpl_m_mdata,
    input  logic                                               i_aic_4_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_aic_5_aon_clk,
    input  wire                                                i_aic_5_aon_rst_n,
    input  wire                                                i_aic_5_clk,
    input  wire                                                i_aic_5_clken,
    input  chip_pkg::chip_axi_addr_t                           i_aic_5_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_5_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_5_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_5_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_5_init_ht_axi_s_arlen,
    input  logic                                               i_aic_5_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_5_init_ht_axi_s_arprot,
    output logic                                               o_aic_5_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_5_init_ht_axi_s_arsize,
    input  logic                                               i_aic_5_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_aic_5_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_5_init_ht_axi_s_rid,
    output logic                                               o_aic_5_init_ht_axi_s_rlast,
    input  logic                                               i_aic_5_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_5_init_ht_axi_s_rresp,
    output logic                                               o_aic_5_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_5_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_5_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_5_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_5_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_5_init_ht_axi_s_awlen,
    input  logic                                               i_aic_5_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_5_init_ht_axi_s_awprot,
    output logic                                               o_aic_5_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_5_init_ht_axi_s_awsize,
    input  logic                                               i_aic_5_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_5_init_ht_axi_s_bid,
    input  logic                                               i_aic_5_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_5_init_ht_axi_s_bresp,
    output logic                                               o_aic_5_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_aic_5_init_ht_axi_s_wdata,
    input  logic                                               i_aic_5_init_ht_axi_s_wlast,
    output logic                                               o_aic_5_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_aic_5_init_ht_axi_s_wstrb,
    input  logic                                               i_aic_5_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_5_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_5_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_5_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_5_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_5_init_lt_axi_s_arlen,
    input  logic                                               i_aic_5_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_5_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_aic_5_init_lt_axi_s_arqos,
    output logic                                               o_aic_5_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_5_init_lt_axi_s_arsize,
    input  logic                                               i_aic_5_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_5_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_5_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_5_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_5_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_5_init_lt_axi_s_awlen,
    input  logic                                               i_aic_5_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_5_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_aic_5_init_lt_axi_s_awqos,
    output logic                                               o_aic_5_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_5_init_lt_axi_s_awsize,
    input  logic                                               i_aic_5_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_5_init_lt_axi_s_bid,
    input  logic                                               i_aic_5_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_5_init_lt_axi_s_bresp,
    output logic                                               o_aic_5_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_5_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_5_init_lt_axi_s_rid,
    output logic                                               o_aic_5_init_lt_axi_s_rlast,
    input  logic                                               i_aic_5_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_5_init_lt_axi_s_rresp,
    output logic                                               o_aic_5_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_5_init_lt_axi_s_wdata,
    input  logic                                               i_aic_5_init_lt_axi_s_wlast,
    output logic                                               o_aic_5_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_aic_5_init_lt_axi_s_wstrb,
    input  logic                                               i_aic_5_init_lt_axi_s_wvalid,
    output logic                                               o_aic_5_pwr_idle_val,
    output logic                                               o_aic_5_pwr_idle_ack,
    input  logic                                               i_aic_5_pwr_idle_req,
    input  wire                                                i_aic_5_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_aic_5_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_aic_5_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_aic_5_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_5_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_aic_5_targ_lt_axi_m_arlen,
    output logic                                               o_aic_5_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_aic_5_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_aic_5_targ_lt_axi_m_arqos,
    input  logic                                               i_aic_5_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_aic_5_targ_lt_axi_m_arsize,
    output logic                                               o_aic_5_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_aic_5_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_aic_5_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_aic_5_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_5_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_aic_5_targ_lt_axi_m_awlen,
    output logic                                               o_aic_5_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_aic_5_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_aic_5_targ_lt_axi_m_awqos,
    input  logic                                               i_aic_5_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_aic_5_targ_lt_axi_m_awsize,
    output logic                                               o_aic_5_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_5_targ_lt_axi_m_bid,
    output logic                                               o_aic_5_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_aic_5_targ_lt_axi_m_bresp,
    input  logic                                               i_aic_5_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_5_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_5_targ_lt_axi_m_rid,
    input  logic                                               i_aic_5_targ_lt_axi_m_rlast,
    output logic                                               o_aic_5_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_aic_5_targ_lt_axi_m_rresp,
    input  logic                                               i_aic_5_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_5_targ_lt_axi_m_wdata,
    output logic                                               o_aic_5_targ_lt_axi_m_wlast,
    input  logic                                               i_aic_5_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_aic_5_targ_lt_axi_m_wstrb,
    output logic                                               o_aic_5_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_aic_5_targ_syscfg_apb_m_paddr,
    output logic                                               o_aic_5_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_aic_5_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_aic_5_targ_syscfg_apb_m_prdata,
    input  logic                                               i_aic_5_targ_syscfg_apb_m_pready,
    output logic                                               o_aic_5_targ_syscfg_apb_m_psel,
    input  logic                                               i_aic_5_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_aic_5_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_aic_5_targ_syscfg_apb_m_pwdata,
    output logic                                               o_aic_5_targ_syscfg_apb_m_pwrite,
    output logic                                               o_aic_5_pwr_tok_idle_val,
    output logic                                               o_aic_5_pwr_tok_idle_ack,
    input  logic                                               i_aic_5_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_aic_5_init_tok_ocpl_s_maddr,
    input  logic                                               i_aic_5_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_aic_5_init_tok_ocpl_s_mdata,
    output logic                                               o_aic_5_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_aic_5_targ_tok_ocpl_m_maddr,
    output logic                                               o_aic_5_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_aic_5_targ_tok_ocpl_m_mdata,
    input  logic                                               i_aic_5_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_aic_6_aon_clk,
    input  wire                                                i_aic_6_aon_rst_n,
    input  wire                                                i_aic_6_clk,
    input  wire                                                i_aic_6_clken,
    input  chip_pkg::chip_axi_addr_t                           i_aic_6_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_6_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_6_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_6_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_6_init_ht_axi_s_arlen,
    input  logic                                               i_aic_6_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_6_init_ht_axi_s_arprot,
    output logic                                               o_aic_6_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_6_init_ht_axi_s_arsize,
    input  logic                                               i_aic_6_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_aic_6_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_6_init_ht_axi_s_rid,
    output logic                                               o_aic_6_init_ht_axi_s_rlast,
    input  logic                                               i_aic_6_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_6_init_ht_axi_s_rresp,
    output logic                                               o_aic_6_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_6_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_6_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_6_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_6_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_6_init_ht_axi_s_awlen,
    input  logic                                               i_aic_6_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_6_init_ht_axi_s_awprot,
    output logic                                               o_aic_6_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_6_init_ht_axi_s_awsize,
    input  logic                                               i_aic_6_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_6_init_ht_axi_s_bid,
    input  logic                                               i_aic_6_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_6_init_ht_axi_s_bresp,
    output logic                                               o_aic_6_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_aic_6_init_ht_axi_s_wdata,
    input  logic                                               i_aic_6_init_ht_axi_s_wlast,
    output logic                                               o_aic_6_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_aic_6_init_ht_axi_s_wstrb,
    input  logic                                               i_aic_6_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_6_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_6_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_6_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_6_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_6_init_lt_axi_s_arlen,
    input  logic                                               i_aic_6_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_6_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_aic_6_init_lt_axi_s_arqos,
    output logic                                               o_aic_6_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_6_init_lt_axi_s_arsize,
    input  logic                                               i_aic_6_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_6_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_6_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_6_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_6_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_6_init_lt_axi_s_awlen,
    input  logic                                               i_aic_6_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_6_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_aic_6_init_lt_axi_s_awqos,
    output logic                                               o_aic_6_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_6_init_lt_axi_s_awsize,
    input  logic                                               i_aic_6_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_6_init_lt_axi_s_bid,
    input  logic                                               i_aic_6_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_6_init_lt_axi_s_bresp,
    output logic                                               o_aic_6_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_6_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_6_init_lt_axi_s_rid,
    output logic                                               o_aic_6_init_lt_axi_s_rlast,
    input  logic                                               i_aic_6_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_6_init_lt_axi_s_rresp,
    output logic                                               o_aic_6_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_6_init_lt_axi_s_wdata,
    input  logic                                               i_aic_6_init_lt_axi_s_wlast,
    output logic                                               o_aic_6_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_aic_6_init_lt_axi_s_wstrb,
    input  logic                                               i_aic_6_init_lt_axi_s_wvalid,
    output logic                                               o_aic_6_pwr_idle_val,
    output logic                                               o_aic_6_pwr_idle_ack,
    input  logic                                               i_aic_6_pwr_idle_req,
    input  wire                                                i_aic_6_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_aic_6_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_aic_6_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_aic_6_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_6_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_aic_6_targ_lt_axi_m_arlen,
    output logic                                               o_aic_6_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_aic_6_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_aic_6_targ_lt_axi_m_arqos,
    input  logic                                               i_aic_6_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_aic_6_targ_lt_axi_m_arsize,
    output logic                                               o_aic_6_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_aic_6_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_aic_6_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_aic_6_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_6_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_aic_6_targ_lt_axi_m_awlen,
    output logic                                               o_aic_6_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_aic_6_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_aic_6_targ_lt_axi_m_awqos,
    input  logic                                               i_aic_6_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_aic_6_targ_lt_axi_m_awsize,
    output logic                                               o_aic_6_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_6_targ_lt_axi_m_bid,
    output logic                                               o_aic_6_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_aic_6_targ_lt_axi_m_bresp,
    input  logic                                               i_aic_6_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_6_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_6_targ_lt_axi_m_rid,
    input  logic                                               i_aic_6_targ_lt_axi_m_rlast,
    output logic                                               o_aic_6_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_aic_6_targ_lt_axi_m_rresp,
    input  logic                                               i_aic_6_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_6_targ_lt_axi_m_wdata,
    output logic                                               o_aic_6_targ_lt_axi_m_wlast,
    input  logic                                               i_aic_6_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_aic_6_targ_lt_axi_m_wstrb,
    output logic                                               o_aic_6_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_aic_6_targ_syscfg_apb_m_paddr,
    output logic                                               o_aic_6_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_aic_6_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_aic_6_targ_syscfg_apb_m_prdata,
    input  logic                                               i_aic_6_targ_syscfg_apb_m_pready,
    output logic                                               o_aic_6_targ_syscfg_apb_m_psel,
    input  logic                                               i_aic_6_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_aic_6_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_aic_6_targ_syscfg_apb_m_pwdata,
    output logic                                               o_aic_6_targ_syscfg_apb_m_pwrite,
    output logic                                               o_aic_6_pwr_tok_idle_val,
    output logic                                               o_aic_6_pwr_tok_idle_ack,
    input  logic                                               i_aic_6_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_aic_6_init_tok_ocpl_s_maddr,
    input  logic                                               i_aic_6_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_aic_6_init_tok_ocpl_s_mdata,
    output logic                                               o_aic_6_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_aic_6_targ_tok_ocpl_m_maddr,
    output logic                                               o_aic_6_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_aic_6_targ_tok_ocpl_m_mdata,
    input  logic                                               i_aic_6_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_aic_7_aon_clk,
    input  wire                                                i_aic_7_aon_rst_n,
    input  wire                                                i_aic_7_clk,
    input  wire                                                i_aic_7_clken,
    input  chip_pkg::chip_axi_addr_t                           i_aic_7_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_7_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_7_init_ht_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_7_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_7_init_ht_axi_s_arlen,
    input  logic                                               i_aic_7_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_7_init_ht_axi_s_arprot,
    output logic                                               o_aic_7_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_7_init_ht_axi_s_arsize,
    input  logic                                               i_aic_7_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_aic_7_init_ht_axi_s_rdata,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_7_init_ht_axi_s_rid,
    output logic                                               o_aic_7_init_ht_axi_s_rlast,
    input  logic                                               i_aic_7_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_7_init_ht_axi_s_rresp,
    output logic                                               o_aic_7_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_7_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_7_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_7_init_ht_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_ht_axi_id_t               i_aic_7_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_7_init_ht_axi_s_awlen,
    input  logic                                               i_aic_7_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_7_init_ht_axi_s_awprot,
    output logic                                               o_aic_7_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_7_init_ht_axi_s_awsize,
    input  logic                                               i_aic_7_init_ht_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_ht_axi_id_t               o_aic_7_init_ht_axi_s_bid,
    input  logic                                               i_aic_7_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_7_init_ht_axi_s_bresp,
    output logic                                               o_aic_7_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_aic_7_init_ht_axi_s_wdata,
    input  logic                                               i_aic_7_init_ht_axi_s_wlast,
    output logic                                               o_aic_7_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_aic_7_init_ht_axi_s_wstrb,
    input  logic                                               i_aic_7_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_7_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_aic_7_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_aic_7_init_lt_axi_s_arcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_7_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_aic_7_init_lt_axi_s_arlen,
    input  logic                                               i_aic_7_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_aic_7_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_aic_7_init_lt_axi_s_arqos,
    output logic                                               o_aic_7_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_aic_7_init_lt_axi_s_arsize,
    input  logic                                               i_aic_7_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_aic_7_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_aic_7_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_aic_7_init_lt_axi_s_awcache,
    input  ai_core_pkg::ai_core_init_lt_axi_id_t               i_aic_7_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_aic_7_init_lt_axi_s_awlen,
    input  logic                                               i_aic_7_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_aic_7_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_aic_7_init_lt_axi_s_awqos,
    output logic                                               o_aic_7_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_aic_7_init_lt_axi_s_awsize,
    input  logic                                               i_aic_7_init_lt_axi_s_awvalid,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_7_init_lt_axi_s_bid,
    input  logic                                               i_aic_7_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_aic_7_init_lt_axi_s_bresp,
    output logic                                               o_aic_7_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_7_init_lt_axi_s_rdata,
    output ai_core_pkg::ai_core_init_lt_axi_id_t               o_aic_7_init_lt_axi_s_rid,
    output logic                                               o_aic_7_init_lt_axi_s_rlast,
    input  logic                                               i_aic_7_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_aic_7_init_lt_axi_s_rresp,
    output logic                                               o_aic_7_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_7_init_lt_axi_s_wdata,
    input  logic                                               i_aic_7_init_lt_axi_s_wlast,
    output logic                                               o_aic_7_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_aic_7_init_lt_axi_s_wstrb,
    input  logic                                               i_aic_7_init_lt_axi_s_wvalid,
    output logic                                               o_aic_7_pwr_idle_val,
    output logic                                               o_aic_7_pwr_idle_ack,
    input  logic                                               i_aic_7_pwr_idle_req,
    input  wire                                                i_aic_7_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_aic_7_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_aic_7_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_aic_7_targ_lt_axi_m_arcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_7_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_aic_7_targ_lt_axi_m_arlen,
    output logic                                               o_aic_7_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_aic_7_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_aic_7_targ_lt_axi_m_arqos,
    input  logic                                               i_aic_7_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_aic_7_targ_lt_axi_m_arsize,
    output logic                                               o_aic_7_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_aic_7_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_aic_7_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_aic_7_targ_lt_axi_m_awcache,
    output ai_core_pkg::ai_core_targ_lt_axi_id_t               o_aic_7_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_aic_7_targ_lt_axi_m_awlen,
    output logic                                               o_aic_7_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_aic_7_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_aic_7_targ_lt_axi_m_awqos,
    input  logic                                               i_aic_7_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_aic_7_targ_lt_axi_m_awsize,
    output logic                                               o_aic_7_targ_lt_axi_m_awvalid,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_7_targ_lt_axi_m_bid,
    output logic                                               o_aic_7_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_aic_7_targ_lt_axi_m_bresp,
    input  logic                                               i_aic_7_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_aic_7_targ_lt_axi_m_rdata,
    input  ai_core_pkg::ai_core_targ_lt_axi_id_t               i_aic_7_targ_lt_axi_m_rid,
    input  logic                                               i_aic_7_targ_lt_axi_m_rlast,
    output logic                                               o_aic_7_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_aic_7_targ_lt_axi_m_rresp,
    input  logic                                               i_aic_7_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_aic_7_targ_lt_axi_m_wdata,
    output logic                                               o_aic_7_targ_lt_axi_m_wlast,
    input  logic                                               i_aic_7_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_aic_7_targ_lt_axi_m_wstrb,
    output logic                                               o_aic_7_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_aic_7_targ_syscfg_apb_m_paddr,
    output logic                                               o_aic_7_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_aic_7_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_aic_7_targ_syscfg_apb_m_prdata,
    input  logic                                               i_aic_7_targ_syscfg_apb_m_pready,
    output logic                                               o_aic_7_targ_syscfg_apb_m_psel,
    input  logic                                               i_aic_7_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_aic_7_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_aic_7_targ_syscfg_apb_m_pwdata,
    output logic                                               o_aic_7_targ_syscfg_apb_m_pwrite,
    output logic                                               o_aic_7_pwr_tok_idle_val,
    output logic                                               o_aic_7_pwr_tok_idle_ack,
    input  logic                                               i_aic_7_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_aic_7_init_tok_ocpl_s_maddr,
    input  logic                                               i_aic_7_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_aic_7_init_tok_ocpl_s_mdata,
    output logic                                               o_aic_7_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_aic_7_targ_tok_ocpl_m_maddr,
    output logic                                               o_aic_7_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_aic_7_targ_tok_ocpl_m_mdata,
    input  logic                                               i_aic_7_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_apu_aon_clk,
    input  wire                                                i_apu_aon_rst_n,
    input  chip_pkg::chip_axi_addr_t                           i_apu_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_apu_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_apu_init_lt_axi_s_arcache,
    input  logic[9:0]                                          i_apu_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_apu_init_lt_axi_s_arlen,
    input  logic                                               i_apu_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_apu_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_apu_init_lt_axi_s_arqos,
    output logic                                               o_apu_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_apu_init_lt_axi_s_arsize,
    input  logic                                               i_apu_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_apu_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_apu_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_apu_init_lt_axi_s_awcache,
    input  logic[9:0]                                          i_apu_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_apu_init_lt_axi_s_awlen,
    input  logic                                               i_apu_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_apu_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_apu_init_lt_axi_s_awqos,
    output logic                                               o_apu_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_apu_init_lt_axi_s_awsize,
    input  logic                                               i_apu_init_lt_axi_s_awvalid,
    output logic[9:0]                                          o_apu_init_lt_axi_s_bid,
    input  logic                                               i_apu_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_apu_init_lt_axi_s_bresp,
    output logic                                               o_apu_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_apu_init_lt_axi_s_rdata,
    output logic[9:0]                                          o_apu_init_lt_axi_s_rid,
    output logic                                               o_apu_init_lt_axi_s_rlast,
    input  logic                                               i_apu_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_apu_init_lt_axi_s_rresp,
    output logic                                               o_apu_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_apu_init_lt_axi_s_wdata,
    input  logic                                               i_apu_init_lt_axi_s_wlast,
    output logic                                               o_apu_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_apu_init_lt_axi_s_wstrb,
    input  logic                                               i_apu_init_lt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_apu_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_apu_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_apu_init_mt_axi_s_arcache,
    input  logic[8:0]                                          i_apu_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_apu_init_mt_axi_s_arlen,
    input  logic                                               i_apu_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_apu_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_apu_init_mt_axi_s_arqos,
    output logic                                               o_apu_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_apu_init_mt_axi_s_arsize,
    input  logic                                               i_apu_init_mt_axi_s_arvalid,
    output apu_pkg::apu_axi_mt_data_t                          o_apu_init_mt_axi_s_rdata,
    output logic[8:0]                                          o_apu_init_mt_axi_s_rid,
    output logic                                               o_apu_init_mt_axi_s_rlast,
    input  logic                                               i_apu_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_apu_init_mt_axi_s_rresp,
    output logic                                               o_apu_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_apu_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_apu_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_apu_init_mt_axi_s_awcache,
    input  logic[8:0]                                          i_apu_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_apu_init_mt_axi_s_awlen,
    input  logic                                               i_apu_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_apu_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_apu_init_mt_axi_s_awqos,
    output logic                                               o_apu_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_apu_init_mt_axi_s_awsize,
    input  logic                                               i_apu_init_mt_axi_s_awvalid,
    output logic[8:0]                                          o_apu_init_mt_axi_s_bid,
    input  logic                                               i_apu_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_apu_init_mt_axi_s_bresp,
    output logic                                               o_apu_init_mt_axi_s_bvalid,
    input  apu_pkg::apu_axi_mt_data_t                          i_apu_init_mt_axi_s_wdata,
    input  logic                                               i_apu_init_mt_axi_s_wlast,
    output logic                                               o_apu_init_mt_axi_s_wready,
    input  apu_pkg::apu_axi_mt_wstrb_t                         i_apu_init_mt_axi_s_wstrb,
    input  logic                                               i_apu_init_mt_axi_s_wvalid,
    output logic                                               o_apu_pwr_idle_val,
    output logic                                               o_apu_pwr_idle_ack,
    input  logic                                               i_apu_pwr_idle_req,
    output chip_pkg::chip_axi_addr_t                           o_apu_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_apu_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_apu_targ_lt_axi_m_arcache,
    output logic[7:0]                                          o_apu_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_apu_targ_lt_axi_m_arlen,
    output logic                                               o_apu_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_apu_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_apu_targ_lt_axi_m_arqos,
    input  logic                                               i_apu_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_apu_targ_lt_axi_m_arsize,
    output logic                                               o_apu_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_apu_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_apu_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_apu_targ_lt_axi_m_awcache,
    output logic[7:0]                                          o_apu_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_apu_targ_lt_axi_m_awlen,
    output logic                                               o_apu_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_apu_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_apu_targ_lt_axi_m_awqos,
    input  logic                                               i_apu_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_apu_targ_lt_axi_m_awsize,
    output logic                                               o_apu_targ_lt_axi_m_awvalid,
    input  logic[7:0]                                          i_apu_targ_lt_axi_m_bid,
    output logic                                               o_apu_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_apu_targ_lt_axi_m_bresp,
    input  logic                                               i_apu_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_apu_targ_lt_axi_m_rdata,
    input  logic[7:0]                                          i_apu_targ_lt_axi_m_rid,
    input  logic                                               i_apu_targ_lt_axi_m_rlast,
    output logic                                               o_apu_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_apu_targ_lt_axi_m_rresp,
    input  logic                                               i_apu_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_apu_targ_lt_axi_m_wdata,
    output logic                                               o_apu_targ_lt_axi_m_wlast,
    input  logic                                               i_apu_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_apu_targ_lt_axi_m_wstrb,
    output logic                                               o_apu_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_apu_targ_syscfg_apb_m_paddr,
    output logic                                               o_apu_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_apu_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_apu_targ_syscfg_apb_m_prdata,
    input  logic                                               i_apu_targ_syscfg_apb_m_pready,
    output logic                                               o_apu_targ_syscfg_apb_m_psel,
    input  logic                                               i_apu_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_apu_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_apu_targ_syscfg_apb_m_pwdata,
    output logic                                               o_apu_targ_syscfg_apb_m_pwrite,
    output logic                                               o_apu_pwr_tok_idle_val,
    output logic                                               o_apu_pwr_tok_idle_ack,
    input  logic                                               i_apu_pwr_tok_idle_req,
    input  chip_pkg::chip_ocpl_token_addr_t                    i_apu_init_tok_ocpl_s_maddr,
    input  logic                                               i_apu_init_tok_ocpl_s_mcmd,
    input  chip_pkg::chip_ocpl_token_data_t                    i_apu_init_tok_ocpl_s_mdata,
    output logic                                               o_apu_init_tok_ocpl_s_scmdaccept,
    output chip_pkg::chip_ocpl_token_addr_t                    o_apu_targ_tok_ocpl_m_maddr,
    output logic                                               o_apu_targ_tok_ocpl_m_mcmd,
    output chip_pkg::chip_ocpl_token_data_t                    o_apu_targ_tok_ocpl_m_mdata,
    input  logic                                               i_apu_targ_tok_ocpl_m_scmdaccept,
    input  wire                                                i_apu_x_clk,
    input  wire                                                i_apu_x_clken,
    input  wire                                                i_apu_x_rst_n,
    input  wire                                                i_dcd_aon_clk,
    input  wire                                                i_dcd_aon_rst_n,
    input  wire                                                i_dcd_codec_clk,
    input  wire                                                i_dcd_codec_clken,
    input  wire                                                i_dcd_codec_rst_n,
    input  chip_pkg::chip_axi_addr_t                           i_dcd_dec_0_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_dcd_dec_0_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_dcd_dec_0_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 i_dcd_dec_0_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_dcd_dec_0_init_mt_axi_s_arlen,
    input  logic                                               i_dcd_dec_0_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_dcd_dec_0_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_dcd_dec_0_init_mt_axi_s_arqos,
    output logic                                               o_dcd_dec_0_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_dcd_dec_0_init_mt_axi_s_arsize,
    input  logic                                               i_dcd_dec_0_init_mt_axi_s_arvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_data_t               o_dcd_dec_0_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 o_dcd_dec_0_init_mt_axi_s_rid,
    output logic                                               o_dcd_dec_0_init_mt_axi_s_rlast,
    input  logic                                               i_dcd_dec_0_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_dcd_dec_0_init_mt_axi_s_rresp,
    output logic                                               o_dcd_dec_0_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_dcd_dec_0_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_dcd_dec_0_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_dcd_dec_0_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 i_dcd_dec_0_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_dcd_dec_0_init_mt_axi_s_awlen,
    input  logic                                               i_dcd_dec_0_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_dcd_dec_0_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_dcd_dec_0_init_mt_axi_s_awqos,
    output logic                                               o_dcd_dec_0_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_dcd_dec_0_init_mt_axi_s_awsize,
    input  logic                                               i_dcd_dec_0_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 o_dcd_dec_0_init_mt_axi_s_bid,
    input  logic                                               i_dcd_dec_0_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_dcd_dec_0_init_mt_axi_s_bresp,
    output logic                                               o_dcd_dec_0_init_mt_axi_s_bvalid,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_data_t               i_dcd_dec_0_init_mt_axi_s_wdata,
    input  logic                                               i_dcd_dec_0_init_mt_axi_s_wlast,
    output logic                                               o_dcd_dec_0_init_mt_axi_s_wready,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_strb_t               i_dcd_dec_0_init_mt_axi_s_wstrb,
    input  logic                                               i_dcd_dec_0_init_mt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_dcd_dec_1_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_dcd_dec_1_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_dcd_dec_1_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 i_dcd_dec_1_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_dcd_dec_1_init_mt_axi_s_arlen,
    input  logic                                               i_dcd_dec_1_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_dcd_dec_1_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_dcd_dec_1_init_mt_axi_s_arqos,
    output logic                                               o_dcd_dec_1_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_dcd_dec_1_init_mt_axi_s_arsize,
    input  logic                                               i_dcd_dec_1_init_mt_axi_s_arvalid,
    output dcd_pkg::dcd_dec_1_init_mt_axi_data_t               o_dcd_dec_1_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 o_dcd_dec_1_init_mt_axi_s_rid,
    output logic                                               o_dcd_dec_1_init_mt_axi_s_rlast,
    input  logic                                               i_dcd_dec_1_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_dcd_dec_1_init_mt_axi_s_rresp,
    output logic                                               o_dcd_dec_1_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_dcd_dec_1_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_dcd_dec_1_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_dcd_dec_1_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 i_dcd_dec_1_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_dcd_dec_1_init_mt_axi_s_awlen,
    input  logic                                               i_dcd_dec_1_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_dcd_dec_1_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_dcd_dec_1_init_mt_axi_s_awqos,
    output logic                                               o_dcd_dec_1_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_dcd_dec_1_init_mt_axi_s_awsize,
    input  logic                                               i_dcd_dec_1_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 o_dcd_dec_1_init_mt_axi_s_bid,
    input  logic                                               i_dcd_dec_1_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_dcd_dec_1_init_mt_axi_s_bresp,
    output logic                                               o_dcd_dec_1_init_mt_axi_s_bvalid,
    input  dcd_pkg::dcd_dec_1_init_mt_axi_data_t               i_dcd_dec_1_init_mt_axi_s_wdata,
    input  logic                                               i_dcd_dec_1_init_mt_axi_s_wlast,
    output logic                                               o_dcd_dec_1_init_mt_axi_s_wready,
    input  dcd_pkg::dcd_dec_1_init_mt_axi_strb_t               i_dcd_dec_1_init_mt_axi_s_wstrb,
    input  logic                                               i_dcd_dec_1_init_mt_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_dcd_dec_2_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_dcd_dec_2_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_dcd_dec_2_init_mt_axi_s_arcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 i_dcd_dec_2_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_dcd_dec_2_init_mt_axi_s_arlen,
    input  logic                                               i_dcd_dec_2_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_dcd_dec_2_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_dcd_dec_2_init_mt_axi_s_arqos,
    output logic                                               o_dcd_dec_2_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_dcd_dec_2_init_mt_axi_s_arsize,
    input  logic                                               i_dcd_dec_2_init_mt_axi_s_arvalid,
    output logic                                       [127:0] o_dcd_dec_2_init_mt_axi_s_rdata,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 o_dcd_dec_2_init_mt_axi_s_rid,
    output logic                                               o_dcd_dec_2_init_mt_axi_s_rlast,
    input  logic                                               i_dcd_dec_2_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_dcd_dec_2_init_mt_axi_s_rresp,
    output logic                                               o_dcd_dec_2_init_mt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_dcd_dec_2_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_dcd_dec_2_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_dcd_dec_2_init_mt_axi_s_awcache,
    input  dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 i_dcd_dec_2_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_dcd_dec_2_init_mt_axi_s_awlen,
    input  logic                                               i_dcd_dec_2_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_dcd_dec_2_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_dcd_dec_2_init_mt_axi_s_awqos,
    output logic                                               o_dcd_dec_2_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_dcd_dec_2_init_mt_axi_s_awsize,
    input  logic                                               i_dcd_dec_2_init_mt_axi_s_awvalid,
    output dcd_pkg::dcd_dec_0_init_mt_axi_id_t                 o_dcd_dec_2_init_mt_axi_s_bid,
    input  logic                                               i_dcd_dec_2_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_dcd_dec_2_init_mt_axi_s_bresp,
    output logic                                               o_dcd_dec_2_init_mt_axi_s_bvalid,
    input  logic                                       [127:0] i_dcd_dec_2_init_mt_axi_s_wdata,
    input  logic                                               i_dcd_dec_2_init_mt_axi_s_wlast,
    output logic                                               o_dcd_dec_2_init_mt_axi_s_wready,
    input  logic                                       [15:0]  i_dcd_dec_2_init_mt_axi_s_wstrb,
    input  logic                                               i_dcd_dec_2_init_mt_axi_s_wvalid,
    input  wire                                                i_dcd_mcu_clk,
    input  wire                                                i_dcd_mcu_clken,
    input  chip_pkg::chip_axi_addr_t                           i_dcd_mcu_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_dcd_mcu_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_dcd_mcu_init_lt_axi_s_arcache,
    input  dcd_pkg::dcd_mcu_init_lt_axi_id_t                   i_dcd_mcu_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_dcd_mcu_init_lt_axi_s_arlen,
    input  logic                                               i_dcd_mcu_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_dcd_mcu_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_dcd_mcu_init_lt_axi_s_arqos,
    output logic                                               o_dcd_mcu_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_dcd_mcu_init_lt_axi_s_arsize,
    input  logic                                               i_dcd_mcu_init_lt_axi_s_arvalid,
    output dcd_pkg::dcd_mcu_init_lt_axi_data_t                 o_dcd_mcu_init_lt_axi_s_rdata,
    output dcd_pkg::dcd_mcu_init_lt_axi_id_t                   o_dcd_mcu_init_lt_axi_s_rid,
    output logic                                               o_dcd_mcu_init_lt_axi_s_rlast,
    input  logic                                               i_dcd_mcu_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_dcd_mcu_init_lt_axi_s_rresp,
    output logic                                               o_dcd_mcu_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_dcd_mcu_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_dcd_mcu_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_dcd_mcu_init_lt_axi_s_awcache,
    input  dcd_pkg::dcd_mcu_init_lt_axi_id_t                   i_dcd_mcu_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_dcd_mcu_init_lt_axi_s_awlen,
    input  logic                                               i_dcd_mcu_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_dcd_mcu_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_dcd_mcu_init_lt_axi_s_awqos,
    output logic                                               o_dcd_mcu_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_dcd_mcu_init_lt_axi_s_awsize,
    input  logic                                               i_dcd_mcu_init_lt_axi_s_awvalid,
    output dcd_pkg::dcd_mcu_init_lt_axi_id_t                   o_dcd_mcu_init_lt_axi_s_bid,
    input  logic                                               i_dcd_mcu_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_dcd_mcu_init_lt_axi_s_bresp,
    output logic                                               o_dcd_mcu_init_lt_axi_s_bvalid,
    input  dcd_pkg::dcd_mcu_init_lt_axi_data_t                 i_dcd_mcu_init_lt_axi_s_wdata,
    input  logic                                               i_dcd_mcu_init_lt_axi_s_wlast,
    output logic                                               o_dcd_mcu_init_lt_axi_s_wready,
    input  dcd_pkg::dcd_mcu_init_lt_axi_strb_t                 i_dcd_mcu_init_lt_axi_s_wstrb,
    input  logic                                               i_dcd_mcu_init_lt_axi_s_wvalid,
    output logic                                               o_dcd_mcu_pwr_idle_val,
    output logic                                               o_dcd_mcu_pwr_idle_ack,
    input  logic                                               i_dcd_mcu_pwr_idle_req,
    input  wire                                                i_dcd_mcu_rst_n,
    output logic                                               o_dcd_pwr_idle_val,
    output logic                                               o_dcd_pwr_idle_ack,
    input  logic                                               i_dcd_pwr_idle_req,
    output dcd_pkg::dcd_targ_cfg_apb_addr_t                    o_dcd_targ_cfg_apb_m_paddr,
    output logic                                               o_dcd_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_dcd_targ_cfg_apb_m_pprot,
    input  dcd_pkg::dcd_targ_cfg_apb_data_t                    i_dcd_targ_cfg_apb_m_prdata,
    input  logic                                               i_dcd_targ_cfg_apb_m_pready,
    output logic                                               o_dcd_targ_cfg_apb_m_psel,
    input  logic                                               i_dcd_targ_cfg_apb_m_pslverr,
    output dcd_pkg::dcd_targ_cfg_apb_strb_t                    o_dcd_targ_cfg_apb_m_pstrb,
    output dcd_pkg::dcd_targ_cfg_apb_data_t                    o_dcd_targ_cfg_apb_m_pwdata,
    output logic                                               o_dcd_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_syscfg_addr_t                        o_dcd_targ_syscfg_apb_m_paddr,
    output logic                                               o_dcd_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_dcd_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_dcd_targ_syscfg_apb_m_prdata,
    input  logic                                               i_dcd_targ_syscfg_apb_m_pready,
    output logic                                               o_dcd_targ_syscfg_apb_m_psel,
    input  logic                                               i_dcd_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_dcd_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_dcd_targ_syscfg_apb_m_pwdata,
    output logic                                               o_dcd_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_ddr_wpll_aon_clk,
    input  wire                                                i_ddr_wpll_aon_rst_n,
    output chip_pkg::chip_syscfg_addr_t                        o_ddr_wpll_targ_syscfg_apb_m_paddr,
    output logic                                               o_ddr_wpll_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_ddr_wpll_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_ddr_wpll_targ_syscfg_apb_m_prdata,
    input  logic                                               i_ddr_wpll_targ_syscfg_apb_m_pready,
    output logic                                               o_ddr_wpll_targ_syscfg_apb_m_psel,
    input  logic                                               i_ddr_wpll_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_ddr_wpll_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_ddr_wpll_targ_syscfg_apb_m_pwdata,
    output logic                                               o_ddr_wpll_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_l2_0_aon_clk,
    input  wire                                                i_l2_0_aon_rst_n,
    input  wire                                                i_l2_0_clk,
    input  wire                                                i_l2_0_clken,
    output logic                                               o_l2_0_pwr_idle_val,
    output logic                                               o_l2_0_pwr_idle_ack,
    input  logic                                               i_l2_0_pwr_idle_req,
    input  wire                                                i_l2_0_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_l2_0_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_l2_0_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_l2_0_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_0_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_l2_0_targ_ht_axi_m_arlen,
    output logic                                               o_l2_0_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_l2_0_targ_ht_axi_m_arprot,
    input  logic                                               i_l2_0_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_l2_0_targ_ht_axi_m_arsize,
    output logic                                               o_l2_0_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_l2_0_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_0_targ_ht_axi_m_rid,
    input  logic                                               i_l2_0_targ_ht_axi_m_rlast,
    output logic                                               o_l2_0_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_l2_0_targ_ht_axi_m_rresp,
    input  logic                                               i_l2_0_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t                           o_l2_0_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_l2_0_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_l2_0_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_0_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_l2_0_targ_ht_axi_m_awlen,
    output logic                                               o_l2_0_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_l2_0_targ_ht_axi_m_awprot,
    input  logic                                               i_l2_0_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_l2_0_targ_ht_axi_m_awsize,
    output logic                                               o_l2_0_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_0_targ_ht_axi_m_bid,
    output logic                                               o_l2_0_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_l2_0_targ_ht_axi_m_bresp,
    input  logic                                               i_l2_0_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_l2_0_targ_ht_axi_m_wdata,
    output logic                                               o_l2_0_targ_ht_axi_m_wlast,
    input  logic                                               i_l2_0_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t                       o_l2_0_targ_ht_axi_m_wstrb,
    output logic                                               o_l2_0_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_l2_0_targ_syscfg_apb_m_paddr,
    output logic                                               o_l2_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_l2_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_l2_0_targ_syscfg_apb_m_prdata,
    input  logic                                               i_l2_0_targ_syscfg_apb_m_pready,
    output logic                                               o_l2_0_targ_syscfg_apb_m_psel,
    input  logic                                               i_l2_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_l2_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_l2_0_targ_syscfg_apb_m_pwdata,
    output logic                                               o_l2_0_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_l2_1_aon_clk,
    input  wire                                                i_l2_1_aon_rst_n,
    input  wire                                                i_l2_1_clk,
    input  wire                                                i_l2_1_clken,
    output logic                                               o_l2_1_pwr_idle_val,
    output logic                                               o_l2_1_pwr_idle_ack,
    input  logic                                               i_l2_1_pwr_idle_req,
    input  wire                                                i_l2_1_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_l2_1_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_l2_1_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_l2_1_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_1_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_l2_1_targ_ht_axi_m_arlen,
    output logic                                               o_l2_1_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_l2_1_targ_ht_axi_m_arprot,
    input  logic                                               i_l2_1_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_l2_1_targ_ht_axi_m_arsize,
    output logic                                               o_l2_1_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_l2_1_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_1_targ_ht_axi_m_rid,
    input  logic                                               i_l2_1_targ_ht_axi_m_rlast,
    output logic                                               o_l2_1_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_l2_1_targ_ht_axi_m_rresp,
    input  logic                                               i_l2_1_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t                           o_l2_1_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_l2_1_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_l2_1_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_1_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_l2_1_targ_ht_axi_m_awlen,
    output logic                                               o_l2_1_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_l2_1_targ_ht_axi_m_awprot,
    input  logic                                               i_l2_1_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_l2_1_targ_ht_axi_m_awsize,
    output logic                                               o_l2_1_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_1_targ_ht_axi_m_bid,
    output logic                                               o_l2_1_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_l2_1_targ_ht_axi_m_bresp,
    input  logic                                               i_l2_1_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_l2_1_targ_ht_axi_m_wdata,
    output logic                                               o_l2_1_targ_ht_axi_m_wlast,
    input  logic                                               i_l2_1_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t                       o_l2_1_targ_ht_axi_m_wstrb,
    output logic                                               o_l2_1_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_l2_1_targ_syscfg_apb_m_paddr,
    output logic                                               o_l2_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_l2_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_l2_1_targ_syscfg_apb_m_prdata,
    input  logic                                               i_l2_1_targ_syscfg_apb_m_pready,
    output logic                                               o_l2_1_targ_syscfg_apb_m_psel,
    input  logic                                               i_l2_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_l2_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_l2_1_targ_syscfg_apb_m_pwdata,
    output logic                                               o_l2_1_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_l2_2_aon_clk,
    input  wire                                                i_l2_2_aon_rst_n,
    input  wire                                                i_l2_2_clk,
    input  wire                                                i_l2_2_clken,
    output logic                                               o_l2_2_pwr_idle_val,
    output logic                                               o_l2_2_pwr_idle_ack,
    input  logic                                               i_l2_2_pwr_idle_req,
    input  wire                                                i_l2_2_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_l2_2_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_l2_2_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_l2_2_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_2_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_l2_2_targ_ht_axi_m_arlen,
    output logic                                               o_l2_2_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_l2_2_targ_ht_axi_m_arprot,
    input  logic                                               i_l2_2_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_l2_2_targ_ht_axi_m_arsize,
    output logic                                               o_l2_2_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_l2_2_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_2_targ_ht_axi_m_rid,
    input  logic                                               i_l2_2_targ_ht_axi_m_rlast,
    output logic                                               o_l2_2_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_l2_2_targ_ht_axi_m_rresp,
    input  logic                                               i_l2_2_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t                           o_l2_2_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_l2_2_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_l2_2_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_2_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_l2_2_targ_ht_axi_m_awlen,
    output logic                                               o_l2_2_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_l2_2_targ_ht_axi_m_awprot,
    input  logic                                               i_l2_2_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_l2_2_targ_ht_axi_m_awsize,
    output logic                                               o_l2_2_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_2_targ_ht_axi_m_bid,
    output logic                                               o_l2_2_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_l2_2_targ_ht_axi_m_bresp,
    input  logic                                               i_l2_2_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_l2_2_targ_ht_axi_m_wdata,
    output logic                                               o_l2_2_targ_ht_axi_m_wlast,
    input  logic                                               i_l2_2_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t                       o_l2_2_targ_ht_axi_m_wstrb,
    output logic                                               o_l2_2_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_l2_2_targ_syscfg_apb_m_paddr,
    output logic                                               o_l2_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_l2_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_l2_2_targ_syscfg_apb_m_prdata,
    input  logic                                               i_l2_2_targ_syscfg_apb_m_pready,
    output logic                                               o_l2_2_targ_syscfg_apb_m_psel,
    input  logic                                               i_l2_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_l2_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_l2_2_targ_syscfg_apb_m_pwdata,
    output logic                                               o_l2_2_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_l2_3_aon_clk,
    input  wire                                                i_l2_3_aon_rst_n,
    input  wire                                                i_l2_3_clk,
    input  wire                                                i_l2_3_clken,
    output logic                                               o_l2_3_pwr_idle_val,
    output logic                                               o_l2_3_pwr_idle_ack,
    input  logic                                               i_l2_3_pwr_idle_req,
    input  wire                                                i_l2_3_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_l2_3_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_l2_3_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_l2_3_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_3_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_l2_3_targ_ht_axi_m_arlen,
    output logic                                               o_l2_3_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_l2_3_targ_ht_axi_m_arprot,
    input  logic                                               i_l2_3_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_l2_3_targ_ht_axi_m_arsize,
    output logic                                               o_l2_3_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_l2_3_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_3_targ_ht_axi_m_rid,
    input  logic                                               i_l2_3_targ_ht_axi_m_rlast,
    output logic                                               o_l2_3_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_l2_3_targ_ht_axi_m_rresp,
    input  logic                                               i_l2_3_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t                           o_l2_3_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_l2_3_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_l2_3_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_3_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_l2_3_targ_ht_axi_m_awlen,
    output logic                                               o_l2_3_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_l2_3_targ_ht_axi_m_awprot,
    input  logic                                               i_l2_3_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_l2_3_targ_ht_axi_m_awsize,
    output logic                                               o_l2_3_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_3_targ_ht_axi_m_bid,
    output logic                                               o_l2_3_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_l2_3_targ_ht_axi_m_bresp,
    input  logic                                               i_l2_3_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_l2_3_targ_ht_axi_m_wdata,
    output logic                                               o_l2_3_targ_ht_axi_m_wlast,
    input  logic                                               i_l2_3_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t                       o_l2_3_targ_ht_axi_m_wstrb,
    output logic                                               o_l2_3_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_l2_3_targ_syscfg_apb_m_paddr,
    output logic                                               o_l2_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_l2_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_l2_3_targ_syscfg_apb_m_prdata,
    input  logic                                               i_l2_3_targ_syscfg_apb_m_pready,
    output logic                                               o_l2_3_targ_syscfg_apb_m_psel,
    input  logic                                               i_l2_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_l2_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_l2_3_targ_syscfg_apb_m_pwdata,
    output logic                                               o_l2_3_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_l2_4_aon_clk,
    input  wire                                                i_l2_4_aon_rst_n,
    input  wire                                                i_l2_4_clk,
    input  wire                                                i_l2_4_clken,
    output logic                                               o_l2_4_pwr_idle_val,
    output logic                                               o_l2_4_pwr_idle_ack,
    input  logic                                               i_l2_4_pwr_idle_req,
    input  wire                                                i_l2_4_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_l2_4_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_l2_4_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_l2_4_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_4_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_l2_4_targ_ht_axi_m_arlen,
    output logic                                               o_l2_4_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_l2_4_targ_ht_axi_m_arprot,
    input  logic                                               i_l2_4_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_l2_4_targ_ht_axi_m_arsize,
    output logic                                               o_l2_4_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_l2_4_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_4_targ_ht_axi_m_rid,
    input  logic                                               i_l2_4_targ_ht_axi_m_rlast,
    output logic                                               o_l2_4_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_l2_4_targ_ht_axi_m_rresp,
    input  logic                                               i_l2_4_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t                           o_l2_4_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_l2_4_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_l2_4_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_4_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_l2_4_targ_ht_axi_m_awlen,
    output logic                                               o_l2_4_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_l2_4_targ_ht_axi_m_awprot,
    input  logic                                               i_l2_4_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_l2_4_targ_ht_axi_m_awsize,
    output logic                                               o_l2_4_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_4_targ_ht_axi_m_bid,
    output logic                                               o_l2_4_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_l2_4_targ_ht_axi_m_bresp,
    input  logic                                               i_l2_4_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_l2_4_targ_ht_axi_m_wdata,
    output logic                                               o_l2_4_targ_ht_axi_m_wlast,
    input  logic                                               i_l2_4_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t                       o_l2_4_targ_ht_axi_m_wstrb,
    output logic                                               o_l2_4_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_l2_4_targ_syscfg_apb_m_paddr,
    output logic                                               o_l2_4_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_l2_4_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_l2_4_targ_syscfg_apb_m_prdata,
    input  logic                                               i_l2_4_targ_syscfg_apb_m_pready,
    output logic                                               o_l2_4_targ_syscfg_apb_m_psel,
    input  logic                                               i_l2_4_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_l2_4_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_l2_4_targ_syscfg_apb_m_pwdata,
    output logic                                               o_l2_4_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_l2_5_aon_clk,
    input  wire                                                i_l2_5_aon_rst_n,
    input  wire                                                i_l2_5_clk,
    input  wire                                                i_l2_5_clken,
    output logic                                               o_l2_5_pwr_idle_val,
    output logic                                               o_l2_5_pwr_idle_ack,
    input  logic                                               i_l2_5_pwr_idle_req,
    input  wire                                                i_l2_5_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_l2_5_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_l2_5_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_l2_5_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_5_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_l2_5_targ_ht_axi_m_arlen,
    output logic                                               o_l2_5_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_l2_5_targ_ht_axi_m_arprot,
    input  logic                                               i_l2_5_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_l2_5_targ_ht_axi_m_arsize,
    output logic                                               o_l2_5_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_l2_5_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_5_targ_ht_axi_m_rid,
    input  logic                                               i_l2_5_targ_ht_axi_m_rlast,
    output logic                                               o_l2_5_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_l2_5_targ_ht_axi_m_rresp,
    input  logic                                               i_l2_5_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t                           o_l2_5_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_l2_5_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_l2_5_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_5_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_l2_5_targ_ht_axi_m_awlen,
    output logic                                               o_l2_5_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_l2_5_targ_ht_axi_m_awprot,
    input  logic                                               i_l2_5_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_l2_5_targ_ht_axi_m_awsize,
    output logic                                               o_l2_5_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_5_targ_ht_axi_m_bid,
    output logic                                               o_l2_5_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_l2_5_targ_ht_axi_m_bresp,
    input  logic                                               i_l2_5_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_l2_5_targ_ht_axi_m_wdata,
    output logic                                               o_l2_5_targ_ht_axi_m_wlast,
    input  logic                                               i_l2_5_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t                       o_l2_5_targ_ht_axi_m_wstrb,
    output logic                                               o_l2_5_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_l2_5_targ_syscfg_apb_m_paddr,
    output logic                                               o_l2_5_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_l2_5_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_l2_5_targ_syscfg_apb_m_prdata,
    input  logic                                               i_l2_5_targ_syscfg_apb_m_pready,
    output logic                                               o_l2_5_targ_syscfg_apb_m_psel,
    input  logic                                               i_l2_5_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_l2_5_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_l2_5_targ_syscfg_apb_m_pwdata,
    output logic                                               o_l2_5_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_l2_6_aon_clk,
    input  wire                                                i_l2_6_aon_rst_n,
    input  wire                                                i_l2_6_clk,
    input  wire                                                i_l2_6_clken,
    output logic                                               o_l2_6_pwr_idle_val,
    output logic                                               o_l2_6_pwr_idle_ack,
    input  logic                                               i_l2_6_pwr_idle_req,
    input  wire                                                i_l2_6_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_l2_6_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_l2_6_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_l2_6_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_6_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_l2_6_targ_ht_axi_m_arlen,
    output logic                                               o_l2_6_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_l2_6_targ_ht_axi_m_arprot,
    input  logic                                               i_l2_6_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_l2_6_targ_ht_axi_m_arsize,
    output logic                                               o_l2_6_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_l2_6_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_6_targ_ht_axi_m_rid,
    input  logic                                               i_l2_6_targ_ht_axi_m_rlast,
    output logic                                               o_l2_6_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_l2_6_targ_ht_axi_m_rresp,
    input  logic                                               i_l2_6_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t                           o_l2_6_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_l2_6_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_l2_6_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_6_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_l2_6_targ_ht_axi_m_awlen,
    output logic                                               o_l2_6_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_l2_6_targ_ht_axi_m_awprot,
    input  logic                                               i_l2_6_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_l2_6_targ_ht_axi_m_awsize,
    output logic                                               o_l2_6_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_6_targ_ht_axi_m_bid,
    output logic                                               o_l2_6_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_l2_6_targ_ht_axi_m_bresp,
    input  logic                                               i_l2_6_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_l2_6_targ_ht_axi_m_wdata,
    output logic                                               o_l2_6_targ_ht_axi_m_wlast,
    input  logic                                               i_l2_6_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t                       o_l2_6_targ_ht_axi_m_wstrb,
    output logic                                               o_l2_6_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_l2_6_targ_syscfg_apb_m_paddr,
    output logic                                               o_l2_6_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_l2_6_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_l2_6_targ_syscfg_apb_m_prdata,
    input  logic                                               i_l2_6_targ_syscfg_apb_m_pready,
    output logic                                               o_l2_6_targ_syscfg_apb_m_psel,
    input  logic                                               i_l2_6_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_l2_6_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_l2_6_targ_syscfg_apb_m_pwdata,
    output logic                                               o_l2_6_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_l2_7_aon_clk,
    input  wire                                                i_l2_7_aon_rst_n,
    input  wire                                                i_l2_7_clk,
    input  wire                                                i_l2_7_clken,
    output logic                                               o_l2_7_pwr_idle_val,
    output logic                                               o_l2_7_pwr_idle_ack,
    input  logic                                               i_l2_7_pwr_idle_req,
    input  wire                                                i_l2_7_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_l2_7_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_l2_7_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_l2_7_targ_ht_axi_m_arcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_7_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_l2_7_targ_ht_axi_m_arlen,
    output logic                                               o_l2_7_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_l2_7_targ_ht_axi_m_arprot,
    input  logic                                               i_l2_7_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_l2_7_targ_ht_axi_m_arsize,
    output logic                                               o_l2_7_targ_ht_axi_m_arvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_l2_7_targ_ht_axi_m_rdata,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_7_targ_ht_axi_m_rid,
    input  logic                                               i_l2_7_targ_ht_axi_m_rlast,
    output logic                                               o_l2_7_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_l2_7_targ_ht_axi_m_rresp,
    input  logic                                               i_l2_7_targ_ht_axi_m_rvalid,
    output chip_pkg::chip_axi_addr_t                           o_l2_7_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_l2_7_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_l2_7_targ_ht_axi_m_awcache,
    output l2_p_pkg::l2_targ_ht_axi_id_t                       o_l2_7_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_l2_7_targ_ht_axi_m_awlen,
    output logic                                               o_l2_7_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_l2_7_targ_ht_axi_m_awprot,
    input  logic                                               i_l2_7_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_l2_7_targ_ht_axi_m_awsize,
    output logic                                               o_l2_7_targ_ht_axi_m_awvalid,
    input  l2_p_pkg::l2_targ_ht_axi_id_t                       i_l2_7_targ_ht_axi_m_bid,
    output logic                                               o_l2_7_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_l2_7_targ_ht_axi_m_bresp,
    input  logic                                               i_l2_7_targ_ht_axi_m_bvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_l2_7_targ_ht_axi_m_wdata,
    output logic                                               o_l2_7_targ_ht_axi_m_wlast,
    input  logic                                               i_l2_7_targ_ht_axi_m_wready,
    output chip_pkg::chip_axi_ht_wstrb_t                       o_l2_7_targ_ht_axi_m_wstrb,
    output logic                                               o_l2_7_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_l2_7_targ_syscfg_apb_m_paddr,
    output logic                                               o_l2_7_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_l2_7_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_l2_7_targ_syscfg_apb_m_prdata,
    input  logic                                               i_l2_7_targ_syscfg_apb_m_pready,
    output logic                                               o_l2_7_targ_syscfg_apb_m_psel,
    input  logic                                               i_l2_7_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_l2_7_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_l2_7_targ_syscfg_apb_m_pwdata,
    output logic                                               o_l2_7_targ_syscfg_apb_m_pwrite,
    input  logic                                               i_l2_addr_mode_port_b0,
    input  logic                                               i_l2_addr_mode_port_b1,
    input  logic                                               i_l2_intr_mode_port_b0,
    input  logic                                               i_l2_intr_mode_port_b1,
    input  wire                                                i_lpddr_graph_0_aon_clk,
    input  wire                                                i_lpddr_graph_0_aon_rst_n,
    input  wire                                                i_lpddr_graph_0_clk,
    input  wire                                                i_lpddr_graph_0_clken,
    output logic[1:0]                                          o_lpddr_graph_0_pwr_idle_vec_val,
    output logic[1:0]                                          o_lpddr_graph_0_pwr_idle_vec_ack,
    input  logic[1:0]                                          i_lpddr_graph_0_pwr_idle_vec_req,
    input  wire                                                i_lpddr_graph_0_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t           o_lpddr_graph_0_targ_cfg_apb_m_paddr,
    output logic                                               o_lpddr_graph_0_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_graph_0_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           i_lpddr_graph_0_targ_cfg_apb_m_prdata,
    input  logic                                               i_lpddr_graph_0_targ_cfg_apb_m_pready,
    output logic                                               o_lpddr_graph_0_targ_cfg_apb_m_psel,
    input  logic                                               i_lpddr_graph_0_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_lpddr_graph_0_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           o_lpddr_graph_0_targ_cfg_apb_m_pwdata,
    output logic                                               o_lpddr_graph_0_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_graph_0_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_lpddr_graph_0_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_lpddr_graph_0_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             o_lpddr_graph_0_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_lpddr_graph_0_targ_ht_axi_m_arlen,
    output logic                                               o_lpddr_graph_0_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_graph_0_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_graph_0_targ_ht_axi_m_arqos,
    input  logic                                               i_lpddr_graph_0_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_lpddr_graph_0_targ_ht_axi_m_arsize,
    output logic                                               o_lpddr_graph_0_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_graph_0_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_lpddr_graph_0_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_lpddr_graph_0_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             o_lpddr_graph_0_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_lpddr_graph_0_targ_ht_axi_m_awlen,
    output logic                                               o_lpddr_graph_0_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_graph_0_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_graph_0_targ_ht_axi_m_awqos,
    input  logic                                               i_lpddr_graph_0_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_lpddr_graph_0_targ_ht_axi_m_awsize,
    output logic                                               o_lpddr_graph_0_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             i_lpddr_graph_0_targ_ht_axi_m_bid,
    output logic                                               o_lpddr_graph_0_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_graph_0_targ_ht_axi_m_bresp,
    input  logic                                               i_lpddr_graph_0_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t           i_lpddr_graph_0_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             i_lpddr_graph_0_targ_ht_axi_m_rid,
    input  logic                                               i_lpddr_graph_0_targ_ht_axi_m_rlast,
    output logic                                               o_lpddr_graph_0_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_graph_0_targ_ht_axi_m_rresp,
    input  logic                                               i_lpddr_graph_0_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t           o_lpddr_graph_0_targ_ht_axi_m_wdata,
    output logic                                               o_lpddr_graph_0_targ_ht_axi_m_wlast,
    input  logic                                               i_lpddr_graph_0_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t           o_lpddr_graph_0_targ_ht_axi_m_wstrb,
    output logic                                               o_lpddr_graph_0_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_lpddr_graph_0_targ_syscfg_apb_m_paddr,
    output logic                                               o_lpddr_graph_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_graph_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_lpddr_graph_0_targ_syscfg_apb_m_prdata,
    input  logic                                               i_lpddr_graph_0_targ_syscfg_apb_m_pready,
    output logic                                               o_lpddr_graph_0_targ_syscfg_apb_m_psel,
    input  logic                                               i_lpddr_graph_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_lpddr_graph_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_lpddr_graph_0_targ_syscfg_apb_m_pwdata,
    output logic                                               o_lpddr_graph_0_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_lpddr_graph_1_aon_clk,
    input  wire                                                i_lpddr_graph_1_aon_rst_n,
    input  wire                                                i_lpddr_graph_1_clk,
    input  wire                                                i_lpddr_graph_1_clken,
    output logic[1:0]                                          o_lpddr_graph_1_pwr_idle_vec_val,
    output logic[1:0]                                          o_lpddr_graph_1_pwr_idle_vec_ack,
    input  logic[1:0]                                          i_lpddr_graph_1_pwr_idle_vec_req,
    input  wire                                                i_lpddr_graph_1_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t           o_lpddr_graph_1_targ_cfg_apb_m_paddr,
    output logic                                               o_lpddr_graph_1_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_graph_1_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           i_lpddr_graph_1_targ_cfg_apb_m_prdata,
    input  logic                                               i_lpddr_graph_1_targ_cfg_apb_m_pready,
    output logic                                               o_lpddr_graph_1_targ_cfg_apb_m_psel,
    input  logic                                               i_lpddr_graph_1_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_lpddr_graph_1_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           o_lpddr_graph_1_targ_cfg_apb_m_pwdata,
    output logic                                               o_lpddr_graph_1_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_graph_1_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_lpddr_graph_1_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_lpddr_graph_1_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             o_lpddr_graph_1_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_lpddr_graph_1_targ_ht_axi_m_arlen,
    output logic                                               o_lpddr_graph_1_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_graph_1_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_graph_1_targ_ht_axi_m_arqos,
    input  logic                                               i_lpddr_graph_1_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_lpddr_graph_1_targ_ht_axi_m_arsize,
    output logic                                               o_lpddr_graph_1_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_graph_1_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_lpddr_graph_1_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_lpddr_graph_1_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             o_lpddr_graph_1_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_lpddr_graph_1_targ_ht_axi_m_awlen,
    output logic                                               o_lpddr_graph_1_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_graph_1_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_graph_1_targ_ht_axi_m_awqos,
    input  logic                                               i_lpddr_graph_1_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_lpddr_graph_1_targ_ht_axi_m_awsize,
    output logic                                               o_lpddr_graph_1_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             i_lpddr_graph_1_targ_ht_axi_m_bid,
    output logic                                               o_lpddr_graph_1_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_graph_1_targ_ht_axi_m_bresp,
    input  logic                                               i_lpddr_graph_1_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t           i_lpddr_graph_1_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             i_lpddr_graph_1_targ_ht_axi_m_rid,
    input  logic                                               i_lpddr_graph_1_targ_ht_axi_m_rlast,
    output logic                                               o_lpddr_graph_1_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_graph_1_targ_ht_axi_m_rresp,
    input  logic                                               i_lpddr_graph_1_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t           o_lpddr_graph_1_targ_ht_axi_m_wdata,
    output logic                                               o_lpddr_graph_1_targ_ht_axi_m_wlast,
    input  logic                                               i_lpddr_graph_1_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t           o_lpddr_graph_1_targ_ht_axi_m_wstrb,
    output logic                                               o_lpddr_graph_1_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_lpddr_graph_1_targ_syscfg_apb_m_paddr,
    output logic                                               o_lpddr_graph_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_graph_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_lpddr_graph_1_targ_syscfg_apb_m_prdata,
    input  logic                                               i_lpddr_graph_1_targ_syscfg_apb_m_pready,
    output logic                                               o_lpddr_graph_1_targ_syscfg_apb_m_psel,
    input  logic                                               i_lpddr_graph_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_lpddr_graph_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_lpddr_graph_1_targ_syscfg_apb_m_pwdata,
    output logic                                               o_lpddr_graph_1_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_lpddr_graph_2_aon_clk,
    input  wire                                                i_lpddr_graph_2_aon_rst_n,
    input  wire                                                i_lpddr_graph_2_clk,
    input  wire                                                i_lpddr_graph_2_clken,
    output logic[1:0]                                          o_lpddr_graph_2_pwr_idle_vec_val,
    output logic[1:0]                                          o_lpddr_graph_2_pwr_idle_vec_ack,
    input  logic[1:0]                                          i_lpddr_graph_2_pwr_idle_vec_req,
    input  wire                                                i_lpddr_graph_2_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t           o_lpddr_graph_2_targ_cfg_apb_m_paddr,
    output logic                                               o_lpddr_graph_2_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_graph_2_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           i_lpddr_graph_2_targ_cfg_apb_m_prdata,
    input  logic                                               i_lpddr_graph_2_targ_cfg_apb_m_pready,
    output logic                                               o_lpddr_graph_2_targ_cfg_apb_m_psel,
    input  logic                                               i_lpddr_graph_2_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_lpddr_graph_2_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           o_lpddr_graph_2_targ_cfg_apb_m_pwdata,
    output logic                                               o_lpddr_graph_2_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_graph_2_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_lpddr_graph_2_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_lpddr_graph_2_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             o_lpddr_graph_2_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_lpddr_graph_2_targ_ht_axi_m_arlen,
    output logic                                               o_lpddr_graph_2_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_graph_2_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_graph_2_targ_ht_axi_m_arqos,
    input  logic                                               i_lpddr_graph_2_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_lpddr_graph_2_targ_ht_axi_m_arsize,
    output logic                                               o_lpddr_graph_2_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_graph_2_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_lpddr_graph_2_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_lpddr_graph_2_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             o_lpddr_graph_2_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_lpddr_graph_2_targ_ht_axi_m_awlen,
    output logic                                               o_lpddr_graph_2_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_graph_2_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_graph_2_targ_ht_axi_m_awqos,
    input  logic                                               i_lpddr_graph_2_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_lpddr_graph_2_targ_ht_axi_m_awsize,
    output logic                                               o_lpddr_graph_2_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             i_lpddr_graph_2_targ_ht_axi_m_bid,
    output logic                                               o_lpddr_graph_2_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_graph_2_targ_ht_axi_m_bresp,
    input  logic                                               i_lpddr_graph_2_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t           i_lpddr_graph_2_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             i_lpddr_graph_2_targ_ht_axi_m_rid,
    input  logic                                               i_lpddr_graph_2_targ_ht_axi_m_rlast,
    output logic                                               o_lpddr_graph_2_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_graph_2_targ_ht_axi_m_rresp,
    input  logic                                               i_lpddr_graph_2_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t           o_lpddr_graph_2_targ_ht_axi_m_wdata,
    output logic                                               o_lpddr_graph_2_targ_ht_axi_m_wlast,
    input  logic                                               i_lpddr_graph_2_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t           o_lpddr_graph_2_targ_ht_axi_m_wstrb,
    output logic                                               o_lpddr_graph_2_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_lpddr_graph_2_targ_syscfg_apb_m_paddr,
    output logic                                               o_lpddr_graph_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_graph_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_lpddr_graph_2_targ_syscfg_apb_m_prdata,
    input  logic                                               i_lpddr_graph_2_targ_syscfg_apb_m_pready,
    output logic                                               o_lpddr_graph_2_targ_syscfg_apb_m_psel,
    input  logic                                               i_lpddr_graph_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_lpddr_graph_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_lpddr_graph_2_targ_syscfg_apb_m_pwdata,
    output logic                                               o_lpddr_graph_2_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_lpddr_graph_3_aon_clk,
    input  wire                                                i_lpddr_graph_3_aon_rst_n,
    input  wire                                                i_lpddr_graph_3_clk,
    input  wire                                                i_lpddr_graph_3_clken,
    output logic[1:0]                                          o_lpddr_graph_3_pwr_idle_vec_val,
    output logic[1:0]                                          o_lpddr_graph_3_pwr_idle_vec_ack,
    input  logic[1:0]                                          i_lpddr_graph_3_pwr_idle_vec_req,
    input  wire                                                i_lpddr_graph_3_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t           o_lpddr_graph_3_targ_cfg_apb_m_paddr,
    output logic                                               o_lpddr_graph_3_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_graph_3_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           i_lpddr_graph_3_targ_cfg_apb_m_prdata,
    input  logic                                               i_lpddr_graph_3_targ_cfg_apb_m_pready,
    output logic                                               o_lpddr_graph_3_targ_cfg_apb_m_psel,
    input  logic                                               i_lpddr_graph_3_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_lpddr_graph_3_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           o_lpddr_graph_3_targ_cfg_apb_m_pwdata,
    output logic                                               o_lpddr_graph_3_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_graph_3_targ_ht_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_lpddr_graph_3_targ_ht_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_lpddr_graph_3_targ_ht_axi_m_arcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             o_lpddr_graph_3_targ_ht_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_lpddr_graph_3_targ_ht_axi_m_arlen,
    output logic                                               o_lpddr_graph_3_targ_ht_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_graph_3_targ_ht_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_graph_3_targ_ht_axi_m_arqos,
    input  logic                                               i_lpddr_graph_3_targ_ht_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_lpddr_graph_3_targ_ht_axi_m_arsize,
    output logic                                               o_lpddr_graph_3_targ_ht_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_graph_3_targ_ht_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_lpddr_graph_3_targ_ht_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_lpddr_graph_3_targ_ht_axi_m_awcache,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             o_lpddr_graph_3_targ_ht_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_lpddr_graph_3_targ_ht_axi_m_awlen,
    output logic                                               o_lpddr_graph_3_targ_ht_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_graph_3_targ_ht_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_graph_3_targ_ht_axi_m_awqos,
    input  logic                                               i_lpddr_graph_3_targ_ht_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_lpddr_graph_3_targ_ht_axi_m_awsize,
    output logic                                               o_lpddr_graph_3_targ_ht_axi_m_awvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             i_lpddr_graph_3_targ_ht_axi_m_bid,
    output logic                                               o_lpddr_graph_3_targ_ht_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_graph_3_targ_ht_axi_m_bresp,
    input  logic                                               i_lpddr_graph_3_targ_ht_axi_m_bvalid,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_data_t           i_lpddr_graph_3_targ_ht_axi_m_rdata,
    input  lpddr_pkg::lpddr_graph_targ_ht_axi_id_t             i_lpddr_graph_3_targ_ht_axi_m_rid,
    input  logic                                               i_lpddr_graph_3_targ_ht_axi_m_rlast,
    output logic                                               o_lpddr_graph_3_targ_ht_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_graph_3_targ_ht_axi_m_rresp,
    input  logic                                               i_lpddr_graph_3_targ_ht_axi_m_rvalid,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_data_t           o_lpddr_graph_3_targ_ht_axi_m_wdata,
    output logic                                               o_lpddr_graph_3_targ_ht_axi_m_wlast,
    input  logic                                               i_lpddr_graph_3_targ_ht_axi_m_wready,
    output lpddr_pkg::lpddr_graph_targ_ht_axi_strb_t           o_lpddr_graph_3_targ_ht_axi_m_wstrb,
    output logic                                               o_lpddr_graph_3_targ_ht_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_lpddr_graph_3_targ_syscfg_apb_m_paddr,
    output logic                                               o_lpddr_graph_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_graph_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_lpddr_graph_3_targ_syscfg_apb_m_prdata,
    input  logic                                               i_lpddr_graph_3_targ_syscfg_apb_m_pready,
    output logic                                               o_lpddr_graph_3_targ_syscfg_apb_m_psel,
    input  logic                                               i_lpddr_graph_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_lpddr_graph_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_lpddr_graph_3_targ_syscfg_apb_m_pwdata,
    output logic                                               o_lpddr_graph_3_targ_syscfg_apb_m_pwrite,
    input  logic                                               i_lpddr_graph_addr_mode_port_b0,
    input  logic                                               i_lpddr_graph_addr_mode_port_b1,
    input  logic                                               i_lpddr_graph_intr_mode_port_b0,
    input  logic                                               i_lpddr_graph_intr_mode_port_b1,
    input  wire                                                i_lpddr_ppp_0_aon_clk,
    input  wire                                                i_lpddr_ppp_0_aon_rst_n,
    input  wire                                                i_lpddr_ppp_0_clk,
    input  wire                                                i_lpddr_ppp_0_clken,
    output logic[1:0]                                          o_lpddr_ppp_0_pwr_idle_vec_val,
    output logic[1:0]                                          o_lpddr_ppp_0_pwr_idle_vec_ack,
    input  logic[1:0]                                          i_lpddr_ppp_0_pwr_idle_vec_req,
    input  wire                                                i_lpddr_ppp_0_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t           o_lpddr_ppp_0_targ_cfg_apb_m_paddr,
    output logic                                               o_lpddr_ppp_0_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_ppp_0_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           i_lpddr_ppp_0_targ_cfg_apb_m_prdata,
    input  logic                                               i_lpddr_ppp_0_targ_cfg_apb_m_pready,
    output logic                                               o_lpddr_ppp_0_targ_cfg_apb_m_psel,
    input  logic                                               i_lpddr_ppp_0_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_lpddr_ppp_0_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           o_lpddr_ppp_0_targ_cfg_apb_m_pwdata,
    output logic                                               o_lpddr_ppp_0_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_ppp_0_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_lpddr_ppp_0_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_lpddr_ppp_0_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               o_lpddr_ppp_0_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_lpddr_ppp_0_targ_mt_axi_m_arlen,
    output logic                                               o_lpddr_ppp_0_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_ppp_0_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_ppp_0_targ_mt_axi_m_arqos,
    input  logic                                               i_lpddr_ppp_0_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_lpddr_ppp_0_targ_mt_axi_m_arsize,
    output logic                                               o_lpddr_ppp_0_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_ppp_0_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_lpddr_ppp_0_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_lpddr_ppp_0_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               o_lpddr_ppp_0_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_lpddr_ppp_0_targ_mt_axi_m_awlen,
    output logic                                               o_lpddr_ppp_0_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_ppp_0_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_ppp_0_targ_mt_axi_m_awqos,
    input  logic                                               i_lpddr_ppp_0_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_lpddr_ppp_0_targ_mt_axi_m_awsize,
    output logic                                               o_lpddr_ppp_0_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               i_lpddr_ppp_0_targ_mt_axi_m_bid,
    output logic                                               o_lpddr_ppp_0_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_ppp_0_targ_mt_axi_m_bresp,
    input  logic                                               i_lpddr_ppp_0_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t             i_lpddr_ppp_0_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               i_lpddr_ppp_0_targ_mt_axi_m_rid,
    input  logic                                               i_lpddr_ppp_0_targ_mt_axi_m_rlast,
    output logic                                               o_lpddr_ppp_0_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_ppp_0_targ_mt_axi_m_rresp,
    input  logic                                               i_lpddr_ppp_0_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t             o_lpddr_ppp_0_targ_mt_axi_m_wdata,
    output logic                                               o_lpddr_ppp_0_targ_mt_axi_m_wlast,
    input  logic                                               i_lpddr_ppp_0_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t             o_lpddr_ppp_0_targ_mt_axi_m_wstrb,
    output logic                                               o_lpddr_ppp_0_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_lpddr_ppp_0_targ_syscfg_apb_m_paddr,
    output logic                                               o_lpddr_ppp_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_ppp_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_lpddr_ppp_0_targ_syscfg_apb_m_prdata,
    input  logic                                               i_lpddr_ppp_0_targ_syscfg_apb_m_pready,
    output logic                                               o_lpddr_ppp_0_targ_syscfg_apb_m_psel,
    input  logic                                               i_lpddr_ppp_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_lpddr_ppp_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_lpddr_ppp_0_targ_syscfg_apb_m_pwdata,
    output logic                                               o_lpddr_ppp_0_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_lpddr_ppp_1_aon_clk,
    input  wire                                                i_lpddr_ppp_1_aon_rst_n,
    input  wire                                                i_lpddr_ppp_1_clk,
    input  wire                                                i_lpddr_ppp_1_clken,
    output logic[1:0]                                          o_lpddr_ppp_1_pwr_idle_vec_val,
    output logic[1:0]                                          o_lpddr_ppp_1_pwr_idle_vec_ack,
    input  logic[1:0]                                          i_lpddr_ppp_1_pwr_idle_vec_req,
    input  wire                                                i_lpddr_ppp_1_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t           o_lpddr_ppp_1_targ_cfg_apb_m_paddr,
    output logic                                               o_lpddr_ppp_1_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_ppp_1_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           i_lpddr_ppp_1_targ_cfg_apb_m_prdata,
    input  logic                                               i_lpddr_ppp_1_targ_cfg_apb_m_pready,
    output logic                                               o_lpddr_ppp_1_targ_cfg_apb_m_psel,
    input  logic                                               i_lpddr_ppp_1_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_lpddr_ppp_1_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           o_lpddr_ppp_1_targ_cfg_apb_m_pwdata,
    output logic                                               o_lpddr_ppp_1_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_ppp_1_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_lpddr_ppp_1_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_lpddr_ppp_1_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               o_lpddr_ppp_1_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_lpddr_ppp_1_targ_mt_axi_m_arlen,
    output logic                                               o_lpddr_ppp_1_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_ppp_1_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_ppp_1_targ_mt_axi_m_arqos,
    input  logic                                               i_lpddr_ppp_1_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_lpddr_ppp_1_targ_mt_axi_m_arsize,
    output logic                                               o_lpddr_ppp_1_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_ppp_1_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_lpddr_ppp_1_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_lpddr_ppp_1_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               o_lpddr_ppp_1_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_lpddr_ppp_1_targ_mt_axi_m_awlen,
    output logic                                               o_lpddr_ppp_1_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_ppp_1_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_ppp_1_targ_mt_axi_m_awqos,
    input  logic                                               i_lpddr_ppp_1_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_lpddr_ppp_1_targ_mt_axi_m_awsize,
    output logic                                               o_lpddr_ppp_1_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               i_lpddr_ppp_1_targ_mt_axi_m_bid,
    output logic                                               o_lpddr_ppp_1_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_ppp_1_targ_mt_axi_m_bresp,
    input  logic                                               i_lpddr_ppp_1_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t             i_lpddr_ppp_1_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               i_lpddr_ppp_1_targ_mt_axi_m_rid,
    input  logic                                               i_lpddr_ppp_1_targ_mt_axi_m_rlast,
    output logic                                               o_lpddr_ppp_1_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_ppp_1_targ_mt_axi_m_rresp,
    input  logic                                               i_lpddr_ppp_1_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t             o_lpddr_ppp_1_targ_mt_axi_m_wdata,
    output logic                                               o_lpddr_ppp_1_targ_mt_axi_m_wlast,
    input  logic                                               i_lpddr_ppp_1_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t             o_lpddr_ppp_1_targ_mt_axi_m_wstrb,
    output logic                                               o_lpddr_ppp_1_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_lpddr_ppp_1_targ_syscfg_apb_m_paddr,
    output logic                                               o_lpddr_ppp_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_ppp_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_lpddr_ppp_1_targ_syscfg_apb_m_prdata,
    input  logic                                               i_lpddr_ppp_1_targ_syscfg_apb_m_pready,
    output logic                                               o_lpddr_ppp_1_targ_syscfg_apb_m_psel,
    input  logic                                               i_lpddr_ppp_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_lpddr_ppp_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_lpddr_ppp_1_targ_syscfg_apb_m_pwdata,
    output logic                                               o_lpddr_ppp_1_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_lpddr_ppp_2_aon_clk,
    input  wire                                                i_lpddr_ppp_2_aon_rst_n,
    input  wire                                                i_lpddr_ppp_2_clk,
    input  wire                                                i_lpddr_ppp_2_clken,
    output logic[1:0]                                          o_lpddr_ppp_2_pwr_idle_vec_val,
    output logic[1:0]                                          o_lpddr_ppp_2_pwr_idle_vec_ack,
    input  logic[1:0]                                          i_lpddr_ppp_2_pwr_idle_vec_req,
    input  wire                                                i_lpddr_ppp_2_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t           o_lpddr_ppp_2_targ_cfg_apb_m_paddr,
    output logic                                               o_lpddr_ppp_2_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_ppp_2_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           i_lpddr_ppp_2_targ_cfg_apb_m_prdata,
    input  logic                                               i_lpddr_ppp_2_targ_cfg_apb_m_pready,
    output logic                                               o_lpddr_ppp_2_targ_cfg_apb_m_psel,
    input  logic                                               i_lpddr_ppp_2_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_lpddr_ppp_2_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           o_lpddr_ppp_2_targ_cfg_apb_m_pwdata,
    output logic                                               o_lpddr_ppp_2_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_ppp_2_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_lpddr_ppp_2_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_lpddr_ppp_2_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               o_lpddr_ppp_2_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_lpddr_ppp_2_targ_mt_axi_m_arlen,
    output logic                                               o_lpddr_ppp_2_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_ppp_2_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_ppp_2_targ_mt_axi_m_arqos,
    input  logic                                               i_lpddr_ppp_2_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_lpddr_ppp_2_targ_mt_axi_m_arsize,
    output logic                                               o_lpddr_ppp_2_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_ppp_2_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_lpddr_ppp_2_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_lpddr_ppp_2_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               o_lpddr_ppp_2_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_lpddr_ppp_2_targ_mt_axi_m_awlen,
    output logic                                               o_lpddr_ppp_2_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_ppp_2_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_ppp_2_targ_mt_axi_m_awqos,
    input  logic                                               i_lpddr_ppp_2_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_lpddr_ppp_2_targ_mt_axi_m_awsize,
    output logic                                               o_lpddr_ppp_2_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               i_lpddr_ppp_2_targ_mt_axi_m_bid,
    output logic                                               o_lpddr_ppp_2_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_ppp_2_targ_mt_axi_m_bresp,
    input  logic                                               i_lpddr_ppp_2_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t             i_lpddr_ppp_2_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               i_lpddr_ppp_2_targ_mt_axi_m_rid,
    input  logic                                               i_lpddr_ppp_2_targ_mt_axi_m_rlast,
    output logic                                               o_lpddr_ppp_2_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_ppp_2_targ_mt_axi_m_rresp,
    input  logic                                               i_lpddr_ppp_2_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t             o_lpddr_ppp_2_targ_mt_axi_m_wdata,
    output logic                                               o_lpddr_ppp_2_targ_mt_axi_m_wlast,
    input  logic                                               i_lpddr_ppp_2_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t             o_lpddr_ppp_2_targ_mt_axi_m_wstrb,
    output logic                                               o_lpddr_ppp_2_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_lpddr_ppp_2_targ_syscfg_apb_m_paddr,
    output logic                                               o_lpddr_ppp_2_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_ppp_2_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_lpddr_ppp_2_targ_syscfg_apb_m_prdata,
    input  logic                                               i_lpddr_ppp_2_targ_syscfg_apb_m_pready,
    output logic                                               o_lpddr_ppp_2_targ_syscfg_apb_m_psel,
    input  logic                                               i_lpddr_ppp_2_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_lpddr_ppp_2_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_lpddr_ppp_2_targ_syscfg_apb_m_pwdata,
    output logic                                               o_lpddr_ppp_2_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_lpddr_ppp_3_aon_clk,
    input  wire                                                i_lpddr_ppp_3_aon_rst_n,
    input  wire                                                i_lpddr_ppp_3_clk,
    input  wire                                                i_lpddr_ppp_3_clken,
    output logic[1:0]                                          o_lpddr_ppp_3_pwr_idle_vec_val,
    output logic[1:0]                                          o_lpddr_ppp_3_pwr_idle_vec_ack,
    input  logic[1:0]                                          i_lpddr_ppp_3_pwr_idle_vec_req,
    input  wire                                                i_lpddr_ppp_3_rst_n,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_addr_t           o_lpddr_ppp_3_targ_cfg_apb_m_paddr,
    output logic                                               o_lpddr_ppp_3_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_ppp_3_targ_cfg_apb_m_pprot,
    input  lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           i_lpddr_ppp_3_targ_cfg_apb_m_prdata,
    input  logic                                               i_lpddr_ppp_3_targ_cfg_apb_m_pready,
    output logic                                               o_lpddr_ppp_3_targ_cfg_apb_m_psel,
    input  logic                                               i_lpddr_ppp_3_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_lpddr_ppp_3_targ_cfg_apb_m_pstrb,
    output lpddr_pkg::lpddr_targ_phy_cfg_apb3_data_t           o_lpddr_ppp_3_targ_cfg_apb_m_pwdata,
    output logic                                               o_lpddr_ppp_3_targ_cfg_apb_m_pwrite,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_ppp_3_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_lpddr_ppp_3_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_lpddr_ppp_3_targ_mt_axi_m_arcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               o_lpddr_ppp_3_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_lpddr_ppp_3_targ_mt_axi_m_arlen,
    output logic                                               o_lpddr_ppp_3_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_ppp_3_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_ppp_3_targ_mt_axi_m_arqos,
    input  logic                                               i_lpddr_ppp_3_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_lpddr_ppp_3_targ_mt_axi_m_arsize,
    output logic                                               o_lpddr_ppp_3_targ_mt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_lpddr_ppp_3_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_lpddr_ppp_3_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_lpddr_ppp_3_targ_mt_axi_m_awcache,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               o_lpddr_ppp_3_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_lpddr_ppp_3_targ_mt_axi_m_awlen,
    output logic                                               o_lpddr_ppp_3_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_lpddr_ppp_3_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_lpddr_ppp_3_targ_mt_axi_m_awqos,
    input  logic                                               i_lpddr_ppp_3_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_lpddr_ppp_3_targ_mt_axi_m_awsize,
    output logic                                               o_lpddr_ppp_3_targ_mt_axi_m_awvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               i_lpddr_ppp_3_targ_mt_axi_m_bid,
    output logic                                               o_lpddr_ppp_3_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_ppp_3_targ_mt_axi_m_bresp,
    input  logic                                               i_lpddr_ppp_3_targ_mt_axi_m_bvalid,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t             i_lpddr_ppp_3_targ_mt_axi_m_rdata,
    input  lpddr_pkg::lpddr_ppp_targ_mt_axi_id_t               i_lpddr_ppp_3_targ_mt_axi_m_rid,
    input  logic                                               i_lpddr_ppp_3_targ_mt_axi_m_rlast,
    output logic                                               o_lpddr_ppp_3_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_lpddr_ppp_3_targ_mt_axi_m_rresp,
    input  logic                                               i_lpddr_ppp_3_targ_mt_axi_m_rvalid,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_data_t             o_lpddr_ppp_3_targ_mt_axi_m_wdata,
    output logic                                               o_lpddr_ppp_3_targ_mt_axi_m_wlast,
    input  logic                                               i_lpddr_ppp_3_targ_mt_axi_m_wready,
    output lpddr_pkg::lpddr_ppp_targ_mt_axi_strb_t             o_lpddr_ppp_3_targ_mt_axi_m_wstrb,
    output logic                                               o_lpddr_ppp_3_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_lpddr_ppp_3_targ_syscfg_apb_m_paddr,
    output logic                                               o_lpddr_ppp_3_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_lpddr_ppp_3_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_lpddr_ppp_3_targ_syscfg_apb_m_prdata,
    input  logic                                               i_lpddr_ppp_3_targ_syscfg_apb_m_pready,
    output logic                                               o_lpddr_ppp_3_targ_syscfg_apb_m_psel,
    input  logic                                               i_lpddr_ppp_3_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_lpddr_ppp_3_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_lpddr_ppp_3_targ_syscfg_apb_m_pwdata,
    output logic                                               o_lpddr_ppp_3_targ_syscfg_apb_m_pwrite,
    input  logic                                               i_lpddr_ppp_addr_mode_port_b0,
    input  logic                                               i_lpddr_ppp_addr_mode_port_b1,
    input  logic                                               i_lpddr_ppp_intr_mode_port_b0,
    input  logic                                               i_lpddr_ppp_intr_mode_port_b1,
    input  wire                                                i_noc_clk,
    input  wire                                                i_noc_rst_n,
    input  wire                                                i_pcie_aon_clk,
    input  wire                                                i_pcie_aon_rst_n,
    input  wire                                                i_pcie_init_mt_clk,
    input  wire                                                i_pcie_init_mt_clken,
    output logic                                               o_pcie_init_mt_pwr_idle_val,
    output logic                                               o_pcie_init_mt_pwr_idle_ack,
    input  logic                                               i_pcie_init_mt_pwr_idle_req,
    input  chip_pkg::chip_axi_addr_t                           i_pcie_init_mt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_pcie_init_mt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_pcie_init_mt_axi_s_arcache,
    input  pcie_pkg::pcie_init_mt_axi_id_t                     i_pcie_init_mt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_pcie_init_mt_axi_s_arlen,
    input  logic                                               i_pcie_init_mt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_pcie_init_mt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_pcie_init_mt_axi_s_arqos,
    output logic                                               o_pcie_init_mt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_pcie_init_mt_axi_s_arsize,
    input  logic                                               i_pcie_init_mt_axi_s_arvalid,
    output pcie_pkg::pcie_init_mt_axi_data_t                   o_pcie_init_mt_axi_s_rdata,
    output pcie_pkg::pcie_init_mt_axi_id_t                     o_pcie_init_mt_axi_s_rid,
    output logic                                               o_pcie_init_mt_axi_s_rlast,
    input  logic                                               i_pcie_init_mt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_pcie_init_mt_axi_s_rresp,
    output logic                                               o_pcie_init_mt_axi_s_rvalid,
    input  wire                                                i_pcie_init_mt_rst_n,
    input  chip_pkg::chip_axi_addr_t                           i_pcie_init_mt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_pcie_init_mt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_pcie_init_mt_axi_s_awcache,
    input  pcie_pkg::pcie_init_mt_axi_id_t                     i_pcie_init_mt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_pcie_init_mt_axi_s_awlen,
    input  logic                                               i_pcie_init_mt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_pcie_init_mt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_pcie_init_mt_axi_s_awqos,
    output logic                                               o_pcie_init_mt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_pcie_init_mt_axi_s_awsize,
    input  logic                                               i_pcie_init_mt_axi_s_awvalid,
    output pcie_pkg::pcie_init_mt_axi_id_t                     o_pcie_init_mt_axi_s_bid,
    input  logic                                               i_pcie_init_mt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_pcie_init_mt_axi_s_bresp,
    output logic                                               o_pcie_init_mt_axi_s_bvalid,
    input  pcie_pkg::pcie_init_mt_axi_data_t                   i_pcie_init_mt_axi_s_wdata,
    input  logic                                               i_pcie_init_mt_axi_s_wlast,
    output logic                                               o_pcie_init_mt_axi_s_wready,
    input  pcie_pkg::pcie_init_mt_axi_strb_t                   i_pcie_init_mt_axi_s_wstrb,
    input  logic                                               i_pcie_init_mt_axi_s_wvalid,
    output pcie_pkg::pcie_targ_cfg_apb3_addr_t                 o_pcie_targ_cfg_apb_m_paddr,
    output logic                                               o_pcie_targ_cfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_pcie_targ_cfg_apb_m_pprot,
    input  pcie_pkg::pcie_targ_cfg_apb3_data_t                 i_pcie_targ_cfg_apb_m_prdata,
    input  logic                                               i_pcie_targ_cfg_apb_m_pready,
    output logic                                               o_pcie_targ_cfg_apb_m_psel,
    input  logic                                               i_pcie_targ_cfg_apb_m_pslverr,
    output logic                                       [3:0]   o_pcie_targ_cfg_apb_m_pstrb,
    output pcie_pkg::pcie_targ_cfg_apb3_data_t                 o_pcie_targ_cfg_apb_m_pwdata,
    output logic                                               o_pcie_targ_cfg_apb_m_pwrite,
    input  wire                                                i_pcie_targ_cfg_clk,
    input  wire                                                i_pcie_targ_cfg_clken,
    output chip_pkg::chip_axi_addr_t                           o_pcie_targ_cfg_dbi_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_pcie_targ_cfg_dbi_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_pcie_targ_cfg_dbi_axi_m_arcache,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_id_t                o_pcie_targ_cfg_dbi_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_pcie_targ_cfg_dbi_axi_m_arlen,
    output logic                                               o_pcie_targ_cfg_dbi_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_pcie_targ_cfg_dbi_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_pcie_targ_cfg_dbi_axi_m_arqos,
    input  logic                                               i_pcie_targ_cfg_dbi_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_pcie_targ_cfg_dbi_axi_m_arsize,
    output logic                                               o_pcie_targ_cfg_dbi_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_pcie_targ_cfg_dbi_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_pcie_targ_cfg_dbi_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_pcie_targ_cfg_dbi_axi_m_awcache,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_id_t                o_pcie_targ_cfg_dbi_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_pcie_targ_cfg_dbi_axi_m_awlen,
    output logic                                               o_pcie_targ_cfg_dbi_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_pcie_targ_cfg_dbi_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_pcie_targ_cfg_dbi_axi_m_awqos,
    input  logic                                               i_pcie_targ_cfg_dbi_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_pcie_targ_cfg_dbi_axi_m_awsize,
    output logic                                               o_pcie_targ_cfg_dbi_axi_m_awvalid,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_id_t                i_pcie_targ_cfg_dbi_axi_m_bid,
    output logic                                               o_pcie_targ_cfg_dbi_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_pcie_targ_cfg_dbi_axi_m_bresp,
    input  logic                                               i_pcie_targ_cfg_dbi_axi_m_bvalid,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_data_t              i_pcie_targ_cfg_dbi_axi_m_rdata,
    input  pcie_pkg::pcie_targ_cfg_dbi_axi_id_t                i_pcie_targ_cfg_dbi_axi_m_rid,
    input  logic                                               i_pcie_targ_cfg_dbi_axi_m_rlast,
    output logic                                               o_pcie_targ_cfg_dbi_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_pcie_targ_cfg_dbi_axi_m_rresp,
    input  logic                                               i_pcie_targ_cfg_dbi_axi_m_rvalid,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_data_t              o_pcie_targ_cfg_dbi_axi_m_wdata,
    output logic                                               o_pcie_targ_cfg_dbi_axi_m_wlast,
    input  logic                                               i_pcie_targ_cfg_dbi_axi_m_wready,
    output pcie_pkg::pcie_targ_cfg_dbi_axi_strb_t              o_pcie_targ_cfg_dbi_axi_m_wstrb,
    output logic                                               o_pcie_targ_cfg_dbi_axi_m_wvalid,
    input  wire                                                i_pcie_targ_cfg_dbi_clk,
    input  wire                                                i_pcie_targ_cfg_dbi_clken,
    output logic                                               o_pcie_targ_cfg_dbi_pwr_idle_val,
    output logic                                               o_pcie_targ_cfg_dbi_pwr_idle_ack,
    input  logic                                               i_pcie_targ_cfg_dbi_pwr_idle_req,
    input  wire                                                i_pcie_targ_cfg_dbi_rst_n,
    output logic                                               o_pcie_targ_cfg_pwr_idle_val,
    output logic                                               o_pcie_targ_cfg_pwr_idle_ack,
    input  logic                                               i_pcie_targ_cfg_pwr_idle_req,
    input  wire                                                i_pcie_targ_cfg_rst_n,
    input  wire                                                i_pcie_targ_mt_clk,
    input  wire                                                i_pcie_targ_mt_clken,
    output logic                                               o_pcie_targ_mt_pwr_idle_val,
    output logic                                               o_pcie_targ_mt_pwr_idle_ack,
    input  logic                                               i_pcie_targ_mt_pwr_idle_req,
    output chip_pkg::chip_axi_addr_t                           o_pcie_targ_mt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_pcie_targ_mt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_pcie_targ_mt_axi_m_arcache,
    output pcie_pkg::pcie_targ_mt_axi_id_t                     o_pcie_targ_mt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_pcie_targ_mt_axi_m_arlen,
    output logic                                               o_pcie_targ_mt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_pcie_targ_mt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_pcie_targ_mt_axi_m_arqos,
    input  logic                                               i_pcie_targ_mt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_pcie_targ_mt_axi_m_arsize,
    output logic                                               o_pcie_targ_mt_axi_m_arvalid,
    input  pcie_pkg::pcie_targ_mt_axi_data_t                   i_pcie_targ_mt_axi_m_rdata,
    input  pcie_pkg::pcie_targ_mt_axi_id_t                     i_pcie_targ_mt_axi_m_rid,
    input  logic                                               i_pcie_targ_mt_axi_m_rlast,
    output logic                                               o_pcie_targ_mt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_pcie_targ_mt_axi_m_rresp,
    input  logic                                               i_pcie_targ_mt_axi_m_rvalid,
    input  wire                                                i_pcie_targ_mt_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_pcie_targ_mt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_pcie_targ_mt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_pcie_targ_mt_axi_m_awcache,
    output pcie_pkg::pcie_targ_mt_axi_id_t                     o_pcie_targ_mt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_pcie_targ_mt_axi_m_awlen,
    output logic                                               o_pcie_targ_mt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_pcie_targ_mt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_pcie_targ_mt_axi_m_awqos,
    input  logic                                               i_pcie_targ_mt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_pcie_targ_mt_axi_m_awsize,
    output logic                                               o_pcie_targ_mt_axi_m_awvalid,
    input  pcie_pkg::pcie_targ_mt_axi_id_t                     i_pcie_targ_mt_axi_m_bid,
    output logic                                               o_pcie_targ_mt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_pcie_targ_mt_axi_m_bresp,
    input  logic                                               i_pcie_targ_mt_axi_m_bvalid,
    output pcie_pkg::pcie_targ_mt_axi_data_t                   o_pcie_targ_mt_axi_m_wdata,
    output logic                                               o_pcie_targ_mt_axi_m_wlast,
    input  logic                                               i_pcie_targ_mt_axi_m_wready,
    output pcie_pkg::pcie_targ_mt_axi_strb_t                   o_pcie_targ_mt_axi_m_wstrb,
    output logic                                               o_pcie_targ_mt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_pcie_targ_syscfg_apb_m_paddr,
    output logic                                               o_pcie_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_pcie_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_pcie_targ_syscfg_apb_m_prdata,
    input  logic                                               i_pcie_targ_syscfg_apb_m_pready,
    output logic                                               o_pcie_targ_syscfg_apb_m_psel,
    input  logic                                               i_pcie_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_pcie_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_pcie_targ_syscfg_apb_m_pwdata,
    output logic                                               o_pcie_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_pve_0_aon_clk,
    input  wire                                                i_pve_0_aon_rst_n,
    input  wire                                                i_pve_0_clk,
    input  wire                                                i_pve_0_clken,
    input  chip_pkg::chip_axi_addr_t                           i_pve_0_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_pve_0_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_pve_0_init_ht_axi_s_arcache,
    input  pve_pkg::pve_ht_axi_m_id_t                          i_pve_0_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_pve_0_init_ht_axi_s_arlen,
    input  logic                                               i_pve_0_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_pve_0_init_ht_axi_s_arprot,
    output logic                                               o_pve_0_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_pve_0_init_ht_axi_s_arsize,
    input  logic                                               i_pve_0_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_pve_0_init_ht_axi_s_rdata,
    output pve_pkg::pve_ht_axi_m_id_t                          o_pve_0_init_ht_axi_s_rid,
    output logic                                               o_pve_0_init_ht_axi_s_rlast,
    input  logic                                               i_pve_0_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_pve_0_init_ht_axi_s_rresp,
    output logic                                               o_pve_0_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_pve_0_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_pve_0_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_pve_0_init_ht_axi_s_awcache,
    input  pve_pkg::pve_ht_axi_m_id_t                          i_pve_0_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_pve_0_init_ht_axi_s_awlen,
    input  logic                                               i_pve_0_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_pve_0_init_ht_axi_s_awprot,
    output logic                                               o_pve_0_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_pve_0_init_ht_axi_s_awsize,
    input  logic                                               i_pve_0_init_ht_axi_s_awvalid,
    output pve_pkg::pve_ht_axi_m_id_t                          o_pve_0_init_ht_axi_s_bid,
    input  logic                                               i_pve_0_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_pve_0_init_ht_axi_s_bresp,
    output logic                                               o_pve_0_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_pve_0_init_ht_axi_s_wdata,
    input  logic                                               i_pve_0_init_ht_axi_s_wlast,
    output logic                                               o_pve_0_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_pve_0_init_ht_axi_s_wstrb,
    input  logic                                               i_pve_0_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_pve_0_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_pve_0_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_pve_0_init_lt_axi_s_arcache,
    input  pve_pkg::pve_lt_axi_m_id_t                          i_pve_0_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_pve_0_init_lt_axi_s_arlen,
    input  logic                                               i_pve_0_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_pve_0_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_pve_0_init_lt_axi_s_arqos,
    output logic                                               o_pve_0_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_pve_0_init_lt_axi_s_arsize,
    input  logic                                               i_pve_0_init_lt_axi_s_arvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_pve_0_init_lt_axi_s_rdata,
    output pve_pkg::pve_lt_axi_m_id_t                          o_pve_0_init_lt_axi_s_rid,
    output logic                                               o_pve_0_init_lt_axi_s_rlast,
    input  logic                                               i_pve_0_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_pve_0_init_lt_axi_s_rresp,
    output logic                                               o_pve_0_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_pve_0_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_pve_0_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_pve_0_init_lt_axi_s_awcache,
    input  pve_pkg::pve_lt_axi_m_id_t                          i_pve_0_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_pve_0_init_lt_axi_s_awlen,
    input  logic                                               i_pve_0_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_pve_0_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_pve_0_init_lt_axi_s_awqos,
    output logic                                               o_pve_0_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_pve_0_init_lt_axi_s_awsize,
    input  logic                                               i_pve_0_init_lt_axi_s_awvalid,
    output pve_pkg::pve_lt_axi_m_id_t                          o_pve_0_init_lt_axi_s_bid,
    input  logic                                               i_pve_0_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_pve_0_init_lt_axi_s_bresp,
    output logic                                               o_pve_0_init_lt_axi_s_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_pve_0_init_lt_axi_s_wdata,
    input  logic                                               i_pve_0_init_lt_axi_s_wlast,
    output logic                                               o_pve_0_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_pve_0_init_lt_axi_s_wstrb,
    input  logic                                               i_pve_0_init_lt_axi_s_wvalid,
    output logic                                               o_pve_0_pwr_idle_val,
    output logic                                               o_pve_0_pwr_idle_ack,
    input  logic                                               i_pve_0_pwr_idle_req,
    input  wire                                                i_pve_0_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_pve_0_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_pve_0_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_pve_0_targ_lt_axi_m_arcache,
    output pve_pkg::pve_lt_axi_s_id_t                          o_pve_0_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_pve_0_targ_lt_axi_m_arlen,
    output logic                                               o_pve_0_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_pve_0_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_pve_0_targ_lt_axi_m_arqos,
    input  logic                                               i_pve_0_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_pve_0_targ_lt_axi_m_arsize,
    output logic                                               o_pve_0_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_pve_0_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_pve_0_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_pve_0_targ_lt_axi_m_awcache,
    output pve_pkg::pve_lt_axi_s_id_t                          o_pve_0_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_pve_0_targ_lt_axi_m_awlen,
    output logic                                               o_pve_0_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_pve_0_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_pve_0_targ_lt_axi_m_awqos,
    input  logic                                               i_pve_0_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_pve_0_targ_lt_axi_m_awsize,
    output logic                                               o_pve_0_targ_lt_axi_m_awvalid,
    input  pve_pkg::pve_lt_axi_s_id_t                          i_pve_0_targ_lt_axi_m_bid,
    output logic                                               o_pve_0_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_pve_0_targ_lt_axi_m_bresp,
    input  logic                                               i_pve_0_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_pve_0_targ_lt_axi_m_rdata,
    input  pve_pkg::pve_lt_axi_s_id_t                          i_pve_0_targ_lt_axi_m_rid,
    input  logic                                               i_pve_0_targ_lt_axi_m_rlast,
    output logic                                               o_pve_0_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_pve_0_targ_lt_axi_m_rresp,
    input  logic                                               i_pve_0_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_pve_0_targ_lt_axi_m_wdata,
    output logic                                               o_pve_0_targ_lt_axi_m_wlast,
    input  logic                                               i_pve_0_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_pve_0_targ_lt_axi_m_wstrb,
    output logic                                               o_pve_0_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_pve_0_targ_syscfg_apb_m_paddr,
    output logic                                               o_pve_0_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_pve_0_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_pve_0_targ_syscfg_apb_m_prdata,
    input  logic                                               i_pve_0_targ_syscfg_apb_m_pready,
    output logic                                               o_pve_0_targ_syscfg_apb_m_psel,
    input  logic                                               i_pve_0_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_pve_0_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_pve_0_targ_syscfg_apb_m_pwdata,
    output logic                                               o_pve_0_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_pve_1_aon_clk,
    input  wire                                                i_pve_1_aon_rst_n,
    input  wire                                                i_pve_1_clk,
    input  wire                                                i_pve_1_clken,
    input  chip_pkg::chip_axi_addr_t                           i_pve_1_init_ht_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_pve_1_init_ht_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_pve_1_init_ht_axi_s_arcache,
    input  pve_pkg::pve_ht_axi_m_id_t                          i_pve_1_init_ht_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_pve_1_init_ht_axi_s_arlen,
    input  logic                                               i_pve_1_init_ht_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_pve_1_init_ht_axi_s_arprot,
    output logic                                               o_pve_1_init_ht_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_pve_1_init_ht_axi_s_arsize,
    input  logic                                               i_pve_1_init_ht_axi_s_arvalid,
    output chip_pkg::chip_axi_ht_data_t                        o_pve_1_init_ht_axi_s_rdata,
    output pve_pkg::pve_ht_axi_m_id_t                          o_pve_1_init_ht_axi_s_rid,
    output logic                                               o_pve_1_init_ht_axi_s_rlast,
    input  logic                                               i_pve_1_init_ht_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_pve_1_init_ht_axi_s_rresp,
    output logic                                               o_pve_1_init_ht_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_pve_1_init_ht_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_pve_1_init_ht_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_pve_1_init_ht_axi_s_awcache,
    input  pve_pkg::pve_ht_axi_m_id_t                          i_pve_1_init_ht_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_pve_1_init_ht_axi_s_awlen,
    input  logic                                               i_pve_1_init_ht_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_pve_1_init_ht_axi_s_awprot,
    output logic                                               o_pve_1_init_ht_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_pve_1_init_ht_axi_s_awsize,
    input  logic                                               i_pve_1_init_ht_axi_s_awvalid,
    output pve_pkg::pve_ht_axi_m_id_t                          o_pve_1_init_ht_axi_s_bid,
    input  logic                                               i_pve_1_init_ht_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_pve_1_init_ht_axi_s_bresp,
    output logic                                               o_pve_1_init_ht_axi_s_bvalid,
    input  chip_pkg::chip_axi_ht_data_t                        i_pve_1_init_ht_axi_s_wdata,
    input  logic                                               i_pve_1_init_ht_axi_s_wlast,
    output logic                                               o_pve_1_init_ht_axi_s_wready,
    input  chip_pkg::chip_axi_ht_wstrb_t                       i_pve_1_init_ht_axi_s_wstrb,
    input  logic                                               i_pve_1_init_ht_axi_s_wvalid,
    input  chip_pkg::chip_axi_addr_t                           i_pve_1_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_pve_1_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_pve_1_init_lt_axi_s_arcache,
    input  pve_pkg::pve_lt_axi_m_id_t                          i_pve_1_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_pve_1_init_lt_axi_s_arlen,
    input  logic                                               i_pve_1_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_pve_1_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_pve_1_init_lt_axi_s_arqos,
    output logic                                               o_pve_1_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_pve_1_init_lt_axi_s_arsize,
    input  logic                                               i_pve_1_init_lt_axi_s_arvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_pve_1_init_lt_axi_s_rdata,
    output pve_pkg::pve_lt_axi_m_id_t                          o_pve_1_init_lt_axi_s_rid,
    output logic                                               o_pve_1_init_lt_axi_s_rlast,
    input  logic                                               i_pve_1_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_pve_1_init_lt_axi_s_rresp,
    output logic                                               o_pve_1_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_addr_t                           i_pve_1_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_pve_1_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_pve_1_init_lt_axi_s_awcache,
    input  pve_pkg::pve_lt_axi_m_id_t                          i_pve_1_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_pve_1_init_lt_axi_s_awlen,
    input  logic                                               i_pve_1_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_pve_1_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_pve_1_init_lt_axi_s_awqos,
    output logic                                               o_pve_1_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_pve_1_init_lt_axi_s_awsize,
    input  logic                                               i_pve_1_init_lt_axi_s_awvalid,
    output pve_pkg::pve_lt_axi_m_id_t                          o_pve_1_init_lt_axi_s_bid,
    input  logic                                               i_pve_1_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_pve_1_init_lt_axi_s_bresp,
    output logic                                               o_pve_1_init_lt_axi_s_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_pve_1_init_lt_axi_s_wdata,
    input  logic                                               i_pve_1_init_lt_axi_s_wlast,
    output logic                                               o_pve_1_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_pve_1_init_lt_axi_s_wstrb,
    input  logic                                               i_pve_1_init_lt_axi_s_wvalid,
    output logic                                               o_pve_1_pwr_idle_val,
    output logic                                               o_pve_1_pwr_idle_ack,
    input  logic                                               i_pve_1_pwr_idle_req,
    input  wire                                                i_pve_1_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_pve_1_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_pve_1_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_pve_1_targ_lt_axi_m_arcache,
    output pve_pkg::pve_lt_axi_s_id_t                          o_pve_1_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_pve_1_targ_lt_axi_m_arlen,
    output logic                                               o_pve_1_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_pve_1_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_pve_1_targ_lt_axi_m_arqos,
    input  logic                                               i_pve_1_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_pve_1_targ_lt_axi_m_arsize,
    output logic                                               o_pve_1_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_pve_1_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_pve_1_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_pve_1_targ_lt_axi_m_awcache,
    output pve_pkg::pve_lt_axi_s_id_t                          o_pve_1_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_pve_1_targ_lt_axi_m_awlen,
    output logic                                               o_pve_1_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_pve_1_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_pve_1_targ_lt_axi_m_awqos,
    input  logic                                               i_pve_1_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_pve_1_targ_lt_axi_m_awsize,
    output logic                                               o_pve_1_targ_lt_axi_m_awvalid,
    input  pve_pkg::pve_lt_axi_s_id_t                          i_pve_1_targ_lt_axi_m_bid,
    output logic                                               o_pve_1_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_pve_1_targ_lt_axi_m_bresp,
    input  logic                                               i_pve_1_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_pve_1_targ_lt_axi_m_rdata,
    input  pve_pkg::pve_lt_axi_s_id_t                          i_pve_1_targ_lt_axi_m_rid,
    input  logic                                               i_pve_1_targ_lt_axi_m_rlast,
    output logic                                               o_pve_1_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_pve_1_targ_lt_axi_m_rresp,
    input  logic                                               i_pve_1_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_pve_1_targ_lt_axi_m_wdata,
    output logic                                               o_pve_1_targ_lt_axi_m_wlast,
    input  logic                                               i_pve_1_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_pve_1_targ_lt_axi_m_wstrb,
    output logic                                               o_pve_1_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_pve_1_targ_syscfg_apb_m_paddr,
    output logic                                               o_pve_1_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_pve_1_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_pve_1_targ_syscfg_apb_m_prdata,
    input  logic                                               i_pve_1_targ_syscfg_apb_m_pready,
    output logic                                               o_pve_1_targ_syscfg_apb_m_psel,
    input  logic                                               i_pve_1_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_pve_1_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_pve_1_targ_syscfg_apb_m_pwdata,
    output logic                                               o_pve_1_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_soc_mgmt_aon_clk,
    input  wire                                                i_soc_mgmt_aon_rst_n,
    input  wire                                                i_soc_mgmt_clk,
    input  wire                                                i_soc_mgmt_clken,
    input  chip_pkg::chip_axi_addr_t                           i_soc_mgmt_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_soc_mgmt_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_soc_mgmt_init_lt_axi_s_arcache,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t                i_soc_mgmt_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_soc_mgmt_init_lt_axi_s_arlen,
    input  logic                                               i_soc_mgmt_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_soc_mgmt_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_soc_mgmt_init_lt_axi_s_arqos,
    output logic                                               o_soc_mgmt_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_soc_mgmt_init_lt_axi_s_arsize,
    input  logic                                               i_soc_mgmt_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_soc_mgmt_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_soc_mgmt_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_soc_mgmt_init_lt_axi_s_awcache,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t                i_soc_mgmt_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_soc_mgmt_init_lt_axi_s_awlen,
    input  logic                                               i_soc_mgmt_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_soc_mgmt_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_soc_mgmt_init_lt_axi_s_awqos,
    output logic                                               o_soc_mgmt_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_soc_mgmt_init_lt_axi_s_awsize,
    input  logic                                               i_soc_mgmt_init_lt_axi_s_awvalid,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t                o_soc_mgmt_init_lt_axi_s_bid,
    input  logic                                               i_soc_mgmt_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_soc_mgmt_init_lt_axi_s_bresp,
    output logic                                               o_soc_mgmt_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_soc_mgmt_init_lt_axi_s_rdata,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_m_id_t                o_soc_mgmt_init_lt_axi_s_rid,
    output logic                                               o_soc_mgmt_init_lt_axi_s_rlast,
    input  logic                                               i_soc_mgmt_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_soc_mgmt_init_lt_axi_s_rresp,
    output logic                                               o_soc_mgmt_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_soc_mgmt_init_lt_axi_s_wdata,
    input  logic                                               i_soc_mgmt_init_lt_axi_s_wlast,
    output logic                                               o_soc_mgmt_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_soc_mgmt_init_lt_axi_s_wstrb,
    input  logic                                               i_soc_mgmt_init_lt_axi_s_wvalid,
    output logic                                               o_soc_mgmt_pwr_idle_val,
    output logic                                               o_soc_mgmt_pwr_idle_ack,
    input  logic                                               i_soc_mgmt_pwr_idle_req,
    input  wire                                                i_soc_mgmt_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_soc_mgmt_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_soc_mgmt_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_soc_mgmt_targ_lt_axi_m_arcache,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t                o_soc_mgmt_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_soc_mgmt_targ_lt_axi_m_arlen,
    output logic                                               o_soc_mgmt_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_soc_mgmt_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_soc_mgmt_targ_lt_axi_m_arqos,
    input  logic                                               i_soc_mgmt_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_soc_mgmt_targ_lt_axi_m_arsize,
    output logic                                               o_soc_mgmt_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_soc_mgmt_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_soc_mgmt_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_soc_mgmt_targ_lt_axi_m_awcache,
    output soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t                o_soc_mgmt_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_soc_mgmt_targ_lt_axi_m_awlen,
    output logic                                               o_soc_mgmt_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_soc_mgmt_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_soc_mgmt_targ_lt_axi_m_awqos,
    input  logic                                               i_soc_mgmt_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_soc_mgmt_targ_lt_axi_m_awsize,
    output logic                                               o_soc_mgmt_targ_lt_axi_m_awvalid,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t                i_soc_mgmt_targ_lt_axi_m_bid,
    output logic                                               o_soc_mgmt_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_soc_mgmt_targ_lt_axi_m_bresp,
    input  logic                                               i_soc_mgmt_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_soc_mgmt_targ_lt_axi_m_rdata,
    input  soc_mgmt_pkg::soc_mgmt_lt_axi_s_id_t                i_soc_mgmt_targ_lt_axi_m_rid,
    input  logic                                               i_soc_mgmt_targ_lt_axi_m_rlast,
    output logic                                               o_soc_mgmt_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_soc_mgmt_targ_lt_axi_m_rresp,
    input  logic                                               i_soc_mgmt_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_soc_mgmt_targ_lt_axi_m_wdata,
    output logic                                               o_soc_mgmt_targ_lt_axi_m_wlast,
    input  logic                                               i_soc_mgmt_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_soc_mgmt_targ_lt_axi_m_wstrb,
    output logic                                               o_soc_mgmt_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_soc_mgmt_syscfg_addr_t               o_soc_mgmt_targ_syscfg_apb_m_paddr,
    output logic                                               o_soc_mgmt_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_soc_mgmt_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_soc_mgmt_targ_syscfg_apb_m_prdata,
    input  logic                                               i_soc_mgmt_targ_syscfg_apb_m_pready,
    output logic                                               o_soc_mgmt_targ_syscfg_apb_m_psel,
    input  logic                                               i_soc_mgmt_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_soc_mgmt_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_soc_mgmt_targ_syscfg_apb_m_pwdata,
    output logic                                               o_soc_mgmt_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_soc_periph_aon_clk,
    input  wire                                                i_soc_periph_aon_rst_n,
    input  wire                                                i_soc_periph_clk,
    input  wire                                                i_soc_periph_clken,
    input  chip_pkg::chip_axi_addr_t                           i_soc_periph_init_lt_axi_s_araddr,
    input  axi_pkg::axi_burst_t                                i_soc_periph_init_lt_axi_s_arburst,
    input  axi_pkg::axi_cache_t                                i_soc_periph_init_lt_axi_s_arcache,
    input  soc_periph_pkg::soc_periph_init_lt_axi_id_t         i_soc_periph_init_lt_axi_s_arid,
    input  axi_pkg::axi_len_t                                  i_soc_periph_init_lt_axi_s_arlen,
    input  logic                                               i_soc_periph_init_lt_axi_s_arlock,
    input  axi_pkg::axi_prot_t                                 i_soc_periph_init_lt_axi_s_arprot,
    input  axi_pkg::axi_qos_t                                  i_soc_periph_init_lt_axi_s_arqos,
    output logic                                               o_soc_periph_init_lt_axi_s_arready,
    input  axi_pkg::axi_size_t                                 i_soc_periph_init_lt_axi_s_arsize,
    input  logic                                               i_soc_periph_init_lt_axi_s_arvalid,
    input  chip_pkg::chip_axi_addr_t                           i_soc_periph_init_lt_axi_s_awaddr,
    input  axi_pkg::axi_burst_t                                i_soc_periph_init_lt_axi_s_awburst,
    input  axi_pkg::axi_cache_t                                i_soc_periph_init_lt_axi_s_awcache,
    input  soc_periph_pkg::soc_periph_init_lt_axi_id_t         i_soc_periph_init_lt_axi_s_awid,
    input  axi_pkg::axi_len_t                                  i_soc_periph_init_lt_axi_s_awlen,
    input  logic                                               i_soc_periph_init_lt_axi_s_awlock,
    input  axi_pkg::axi_prot_t                                 i_soc_periph_init_lt_axi_s_awprot,
    input  axi_pkg::axi_qos_t                                  i_soc_periph_init_lt_axi_s_awqos,
    output logic                                               o_soc_periph_init_lt_axi_s_awready,
    input  axi_pkg::axi_size_t                                 i_soc_periph_init_lt_axi_s_awsize,
    input  logic                                               i_soc_periph_init_lt_axi_s_awvalid,
    output soc_periph_pkg::soc_periph_init_lt_axi_id_t         o_soc_periph_init_lt_axi_s_bid,
    input  logic                                               i_soc_periph_init_lt_axi_s_bready,
    output axi_pkg::axi_resp_t                                 o_soc_periph_init_lt_axi_s_bresp,
    output logic                                               o_soc_periph_init_lt_axi_s_bvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_soc_periph_init_lt_axi_s_rdata,
    output soc_periph_pkg::soc_periph_init_lt_axi_id_t         o_soc_periph_init_lt_axi_s_rid,
    output logic                                               o_soc_periph_init_lt_axi_s_rlast,
    input  logic                                               i_soc_periph_init_lt_axi_s_rready,
    output axi_pkg::axi_resp_t                                 o_soc_periph_init_lt_axi_s_rresp,
    output logic                                               o_soc_periph_init_lt_axi_s_rvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_soc_periph_init_lt_axi_s_wdata,
    input  logic                                               i_soc_periph_init_lt_axi_s_wlast,
    output logic                                               o_soc_periph_init_lt_axi_s_wready,
    input  chip_pkg::chip_axi_lt_wstrb_t                       i_soc_periph_init_lt_axi_s_wstrb,
    input  logic                                               i_soc_periph_init_lt_axi_s_wvalid,
    output logic                                               o_soc_periph_pwr_idle_val,
    output logic                                               o_soc_periph_pwr_idle_ack,
    input  logic                                               i_soc_periph_pwr_idle_req,
    input  wire                                                i_soc_periph_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_soc_periph_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_soc_periph_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_soc_periph_targ_lt_axi_m_arcache,
    output soc_periph_pkg::soc_periph_targ_lt_axi_id_t         o_soc_periph_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_soc_periph_targ_lt_axi_m_arlen,
    output logic                                               o_soc_periph_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_soc_periph_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_soc_periph_targ_lt_axi_m_arqos,
    input  logic                                               i_soc_periph_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_soc_periph_targ_lt_axi_m_arsize,
    output logic                                               o_soc_periph_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_soc_periph_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_soc_periph_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_soc_periph_targ_lt_axi_m_awcache,
    output soc_periph_pkg::soc_periph_targ_lt_axi_id_t         o_soc_periph_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_soc_periph_targ_lt_axi_m_awlen,
    output logic                                               o_soc_periph_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_soc_periph_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_soc_periph_targ_lt_axi_m_awqos,
    input  logic                                               i_soc_periph_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_soc_periph_targ_lt_axi_m_awsize,
    output logic                                               o_soc_periph_targ_lt_axi_m_awvalid,
    input  soc_periph_pkg::soc_periph_targ_lt_axi_id_t         i_soc_periph_targ_lt_axi_m_bid,
    output logic                                               o_soc_periph_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_soc_periph_targ_lt_axi_m_bresp,
    input  logic                                               i_soc_periph_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_soc_periph_targ_lt_axi_m_rdata,
    input  soc_periph_pkg::soc_periph_targ_lt_axi_id_t         i_soc_periph_targ_lt_axi_m_rid,
    input  logic                                               i_soc_periph_targ_lt_axi_m_rlast,
    output logic                                               o_soc_periph_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_soc_periph_targ_lt_axi_m_rresp,
    input  logic                                               i_soc_periph_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_soc_periph_targ_lt_axi_m_wdata,
    output logic                                               o_soc_periph_targ_lt_axi_m_wlast,
    input  logic                                               i_soc_periph_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_soc_periph_targ_lt_axi_m_wstrb,
    output logic                                               o_soc_periph_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_soc_periph_targ_syscfg_apb_m_paddr,
    output logic                                               o_soc_periph_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_soc_periph_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_soc_periph_targ_syscfg_apb_m_prdata,
    input  logic                                               i_soc_periph_targ_syscfg_apb_m_pready,
    output logic                                               o_soc_periph_targ_syscfg_apb_m_psel,
    input  logic                                               i_soc_periph_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_soc_periph_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_soc_periph_targ_syscfg_apb_m_pwdata,
    output logic                                               o_soc_periph_targ_syscfg_apb_m_pwrite,
    input  wire                                                i_sys_spm_aon_clk,
    input  wire                                                i_sys_spm_aon_rst_n,
    input  wire                                                i_sys_spm_clk,
    input  wire                                                i_sys_spm_clken,
    output logic                                               o_sys_spm_pwr_idle_val,
    output logic                                               o_sys_spm_pwr_idle_ack,
    input  logic                                               i_sys_spm_pwr_idle_req,
    input  wire                                                i_sys_spm_rst_n,
    output chip_pkg::chip_axi_addr_t                           o_sys_spm_targ_lt_axi_m_araddr,
    output axi_pkg::axi_burst_t                                o_sys_spm_targ_lt_axi_m_arburst,
    output axi_pkg::axi_cache_t                                o_sys_spm_targ_lt_axi_m_arcache,
    output sys_spm_pkg::sys_spm_targ_lt_axi_id_t               o_sys_spm_targ_lt_axi_m_arid,
    output axi_pkg::axi_len_t                                  o_sys_spm_targ_lt_axi_m_arlen,
    output logic                                               o_sys_spm_targ_lt_axi_m_arlock,
    output axi_pkg::axi_prot_t                                 o_sys_spm_targ_lt_axi_m_arprot,
    output axi_pkg::axi_qos_t                                  o_sys_spm_targ_lt_axi_m_arqos,
    input  logic                                               i_sys_spm_targ_lt_axi_m_arready,
    output axi_pkg::axi_size_t                                 o_sys_spm_targ_lt_axi_m_arsize,
    output logic                                               o_sys_spm_targ_lt_axi_m_arvalid,
    output chip_pkg::chip_axi_addr_t                           o_sys_spm_targ_lt_axi_m_awaddr,
    output axi_pkg::axi_burst_t                                o_sys_spm_targ_lt_axi_m_awburst,
    output axi_pkg::axi_cache_t                                o_sys_spm_targ_lt_axi_m_awcache,
    output sys_spm_pkg::sys_spm_targ_lt_axi_id_t               o_sys_spm_targ_lt_axi_m_awid,
    output axi_pkg::axi_len_t                                  o_sys_spm_targ_lt_axi_m_awlen,
    output logic                                               o_sys_spm_targ_lt_axi_m_awlock,
    output axi_pkg::axi_prot_t                                 o_sys_spm_targ_lt_axi_m_awprot,
    output axi_pkg::axi_qos_t                                  o_sys_spm_targ_lt_axi_m_awqos,
    input  logic                                               i_sys_spm_targ_lt_axi_m_awready,
    output axi_pkg::axi_size_t                                 o_sys_spm_targ_lt_axi_m_awsize,
    output logic                                               o_sys_spm_targ_lt_axi_m_awvalid,
    input  sys_spm_pkg::sys_spm_targ_lt_axi_id_t               i_sys_spm_targ_lt_axi_m_bid,
    output logic                                               o_sys_spm_targ_lt_axi_m_bready,
    input  axi_pkg::axi_resp_t                                 i_sys_spm_targ_lt_axi_m_bresp,
    input  logic                                               i_sys_spm_targ_lt_axi_m_bvalid,
    input  chip_pkg::chip_axi_lt_data_t                        i_sys_spm_targ_lt_axi_m_rdata,
    input  sys_spm_pkg::sys_spm_targ_lt_axi_id_t               i_sys_spm_targ_lt_axi_m_rid,
    input  logic                                               i_sys_spm_targ_lt_axi_m_rlast,
    output logic                                               o_sys_spm_targ_lt_axi_m_rready,
    input  axi_pkg::axi_resp_t                                 i_sys_spm_targ_lt_axi_m_rresp,
    input  logic                                               i_sys_spm_targ_lt_axi_m_rvalid,
    output chip_pkg::chip_axi_lt_data_t                        o_sys_spm_targ_lt_axi_m_wdata,
    output logic                                               o_sys_spm_targ_lt_axi_m_wlast,
    input  logic                                               i_sys_spm_targ_lt_axi_m_wready,
    output chip_pkg::chip_axi_lt_wstrb_t                       o_sys_spm_targ_lt_axi_m_wstrb,
    output logic                                               o_sys_spm_targ_lt_axi_m_wvalid,
    output chip_pkg::chip_syscfg_addr_t                        o_sys_spm_targ_syscfg_apb_m_paddr,
    output logic                                               o_sys_spm_targ_syscfg_apb_m_penable,
    output axe_apb_pkg::apb_prot_t                             o_sys_spm_targ_syscfg_apb_m_pprot,
    input  chip_pkg::chip_apb_syscfg_data_t                    i_sys_spm_targ_syscfg_apb_m_prdata,
    input  logic                                               i_sys_spm_targ_syscfg_apb_m_pready,
    output logic                                               o_sys_spm_targ_syscfg_apb_m_psel,
    input  logic                                               i_sys_spm_targ_syscfg_apb_m_pslverr,
    output chip_pkg::chip_apb_syscfg_strb_t                    o_sys_spm_targ_syscfg_apb_m_pstrb,
    output chip_pkg::chip_apb_syscfg_data_t                    o_sys_spm_targ_syscfg_apb_m_pwdata,
    output logic                                               o_sys_spm_targ_syscfg_apb_m_pwrite
);

    // Wire Connections (between subpartitions)
    logic [182:0] dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data;
    logic         dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head;
    logic         dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy;
    logic         dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail;
    logic         dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data;
    logic         dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head;
    logic         dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy;
    logic         dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail;
    logic         dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld;
    logic [398:0] dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data;
    logic         dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head;
    logic         dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld;
    logic [398:0] dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data;
    logic         dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head;
    logic         dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld;
    logic [398:0] dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data;
    logic         dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head;
    logic         dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld;
    logic [398:0] dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data;
    logic         dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head;
    logic         dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld;
    logic [398:0] dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data;
    logic         dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head;
    logic         dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld;
    logic [398:0] dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data;
    logic         dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head;
    logic         dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld;
    logic [398:0] dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data;
    logic         dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head;
    logic         dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld;
    logic [398:0] dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data;
    logic         dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head;
    logic         dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld;
    logic [182:0] dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data;
    logic         dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head;
    logic         dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data;
    logic         dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head;
    logic         dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail;
    logic         dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld;
    logic [398:0] dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data;
    logic         dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head;
    logic         dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy;
    logic         dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail;
    logic         dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld;
    logic [398:0] dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data;
    logic         dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head;
    logic         dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy;
    logic         dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail;
    logic         dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld;
    logic [398:0] dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data;
    logic         dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head;
    logic         dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy;
    logic         dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail;
    logic         dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld;
    logic [398:0] dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data;
    logic         dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head;
    logic         dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy;
    logic         dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail;
    logic         dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld;
    logic [398:0] dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data;
    logic         dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head;
    logic         dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy;
    logic         dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail;
    logic         dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld;
    logic [398:0] dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data;
    logic         dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head;
    logic         dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy;
    logic         dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail;
    logic         dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld;
    logic [398:0] dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data;
    logic         dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head;
    logic         dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy;
    logic         dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail;
    logic         dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld;
    logic [398:0] dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data;
    logic         dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head;
    logic         dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy;
    logic         dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail;
    logic         dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld;
    logic [146:0] dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data;
    logic         dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head;
    logic         dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy;
    logic         dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail;
    logic         dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld;
    logic [146:0] dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data;
    logic         dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head;
    logic         dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy;
    logic         dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail;
    logic         dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld;
    logic [182:0] dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data;
    logic         dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head;
    logic         dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy;
    logic         dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail;
    logic         dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data;
    logic         dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head;
    logic         dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy;
    logic         dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail;
    logic         dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld;
    logic [686:0] dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data;
    logic         dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head;
    logic         dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy;
    logic         dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail;
    logic         dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data;
    logic         dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head;
    logic         dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy;
    logic         dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail;
    logic         dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld;
    logic [686:0] dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data;
    logic         dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head;
    logic         dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy;
    logic         dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail;
    logic         dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data;
    logic         dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head;
    logic         dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy;
    logic         dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail;
    logic         dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld;
    logic [686:0] dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data;
    logic         dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head;
    logic         dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy;
    logic         dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail;
    logic         dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data;
    logic         dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head;
    logic         dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy;
    logic         dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail;
    logic         dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld;
    logic [686:0] dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data;
    logic         dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head;
    logic         dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy;
    logic         dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail;
    logic         dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld;
    logic [182:0] dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data;
    logic         dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head;
    logic         dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy;
    logic         dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail;
    logic         dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld;
    logic [686:0] dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld;
    logic [182:0] dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data;
    logic         dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head;
    logic         dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy;
    logic         dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail;
    logic         dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data;
    logic         dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head;
    logic         dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail;
    logic         dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld;
    logic [686:0] dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data;
    logic         dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head;
    logic         dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy;
    logic         dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail;
    logic         dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data;
    logic         dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head;
    logic         dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data;
    logic         dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head;
    logic         dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy;
    logic         dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail;
    logic         dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data;
    logic         dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head;
    logic         dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld;
    logic [182:0] dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data;
    logic         dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head;
    logic         dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy;
    logic         dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail;
    logic         dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data;
    logic         dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head;
    logic         dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail;
    logic         dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld;
    logic [686:0] dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data;
    logic         dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head;
    logic         dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy;
    logic         dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail;
    logic         dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data;
    logic         dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head;
    logic         dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data;
    logic         dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head;
    logic         dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy;
    logic         dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail;
    logic         dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data;
    logic         dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head;
    logic         dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data;
    logic         dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head;
    logic         dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy;
    logic         dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail;
    logic         dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data;
    logic         dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head;
    logic         dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data;
    logic         dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head;
    logic         dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy;
    logic         dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail;
    logic         dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data;
    logic         dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head;
    logic         dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld;
    logic [182:0] dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data;
    logic         dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head;
    logic         dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy;
    logic         dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail;
    logic         dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data;
    logic         dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head;
    logic         dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail;
    logic         dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld;
    logic [686:0] dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data;
    logic         dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head;
    logic         dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy;
    logic         dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail;
    logic         dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data;
    logic         dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head;
    logic         dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data;
    logic         dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head;
    logic         dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy;
    logic         dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail;
    logic         dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data;
    logic         dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head;
    logic         dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld;
    logic [182:0] dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data;
    logic         dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head;
    logic         dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy;
    logic         dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail;
    logic         dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data;
    logic         dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head;
    logic         dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail;
    logic         dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld;
    logic [182:0] dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data;
    logic         dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head;
    logic         dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy;
    logic         dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail;
    logic         dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data;
    logic         dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head;
    logic         dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail;
    logic         dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data;
    logic         dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head;
    logic         dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail;
    logic         dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data;
    logic         dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head;
    logic         dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail;
    logic         dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data;
    logic         dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head;
    logic         dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail;
    logic         dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data;
    logic         dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head;
    logic         dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail;
    logic         dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data;
    logic         dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head;
    logic         dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail;
    logic         dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data;
    logic         dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head;
    logic         dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail;
    logic         dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data;
    logic         dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head;
    logic         dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail;
    logic         dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data;
    logic         dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head;
    logic         dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail;
    logic         dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data;
    logic         dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head;
    logic         dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail;
    logic         dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data;
    logic         dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head;
    logic         dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail;
    logic         dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data;
    logic         dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head;
    logic         dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail;
    logic         dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data;
    logic         dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head;
    logic         dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy;
    logic         dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail;
    logic         dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data;
    logic         dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head;
    logic         dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld;
    logic [182:0] dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data;
    logic         dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head;
    logic         dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy;
    logic         dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail;
    logic         dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data;
    logic         dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head;
    logic         dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail;
    logic         dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data;
    logic         dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head;
    logic         dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail;
    logic         dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data;
    logic         dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head;
    logic         dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy;
    logic         dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail;
    logic         dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data;
    logic         dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head;
    logic         dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld;
    logic [182:0] dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data;
    logic         dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head;
    logic         dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy;
    logic         dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail;
    logic         dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data;
    logic         dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head;
    logic         dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail;
    logic         dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld;
    logic [146:0] dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data;
    logic         dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head;
    logic         dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail;
    logic         dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data;
    logic         dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head;
    logic         dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail;
    logic         dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data;
    logic         dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head;
    logic         dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail;
    logic         dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data;
    logic         dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head;
    logic         dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail;
    logic         dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data;
    logic         dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head;
    logic         dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail;
    logic         dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data;
    logic         dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head;
    logic         dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail;
    logic         dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data;
    logic         dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head;
    logic         dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail;
    logic         dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data;
    logic         dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head;
    logic         dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail;
    logic         dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data;
    logic         dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head;
    logic         dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail;
    logic         dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld;
    logic [146:0] dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data;
    logic         dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head;
    logic         dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail;
    logic         dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data;
    logic         dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head;
    logic         dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail;
    logic         dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld;
    logic [108:0] dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld;
    logic [146:0] dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data;
    logic         dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head;
    logic         dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy;
    logic         dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail;
    logic         dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld;
    logic [686:0] dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data;
    logic         dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head;
    logic         dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld;
    logic [182:0] dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data;
    logic         dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head;
    logic         dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy;
    logic         dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail;
    logic         dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld;
    logic [182:0] dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data;
    logic         dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head;
    logic         dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy;
    logic         dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail;
    logic         dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld;

    logic [41:0]  dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data;
    logic         dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head;
    logic         dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy;
    logic         dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail;
    logic         dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld;
    logic [31:0]  dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data;
    logic         dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head;
    logic         dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy;
    logic         dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail;
    logic         dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld;
    logic [41:0]  dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data;
    logic         dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head;
    logic         dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy;
    logic         dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail;
    logic         dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld;
    logic [31:0]  dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data;
    logic         dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head;
    logic         dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy;
    logic         dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail;
    logic         dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld;
    logic [41:0]  dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data;
    logic         dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head;
    logic         dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy;
    logic         dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail;
    logic         dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld;
    logic [31:0]  dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data;
    logic         dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head;
    logic         dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy;
    logic         dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail;
    logic         dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld;
    logic [41:0]  dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data;
    logic         dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head;
    logic         dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy;
    logic         dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail;
    logic         dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld;
    logic [31:0]  dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data;
    logic         dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head;
    logic         dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy;
    logic         dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail;
    logic         dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld;
    logic [41:0]  dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data;
    logic         dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head;
    logic         dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy;
    logic         dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail;
    logic         dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld;
    logic [31:0]  dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data;
    logic         dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head;
    logic         dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy;
    logic         dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail;
    logic         dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld;
    logic [41:0]  dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data;
    logic         dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head;
    logic         dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy;
    logic         dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail;
    logic         dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld;
    logic [31:0]  dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data;
    logic         dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head;
    logic         dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy;
    logic         dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail;
    logic         dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld;
    logic [31:0]  dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data;
    logic         dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head;
    logic         dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy;
    logic         dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail;
    logic         dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld;
    logic [41:0]  dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data;
    logic         dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head;
    logic         dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy;
    logic         dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail;
    logic         dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld;
    logic [41:0]  dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data;
    logic         dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head;
    logic         dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy;
    logic         dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail;
    logic         dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld;
    logic [31:0]  dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data;
    logic         dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head;
    logic         dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy;
    logic         dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail;
    logic         dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld;

    // Instance of noc_ddr_east_p
    noc_ddr_east_p ddr_east_p (
        .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data),
        .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head),
        .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy),
        .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail),
        .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld),
        .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data),
        .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head),
        .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy),
        .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail),
        .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data),
        .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head),
        .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data),
        .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head),
        .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld),
        .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
        .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
        .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
        .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
        .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
        .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
        .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
        .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
        .i_lpddr_ppp_0_aon_clk(i_lpddr_ppp_0_aon_clk),
        .i_lpddr_ppp_0_aon_rst_n(i_lpddr_ppp_0_aon_rst_n),
        .o_lpddr_ppp_0_cfg_pwr_idle_val(o_lpddr_ppp_0_pwr_idle_vec_val[0]),
        .o_lpddr_ppp_0_cfg_pwr_idle_ack(o_lpddr_ppp_0_pwr_idle_vec_ack[0]),
        .i_lpddr_ppp_0_cfg_pwr_idle_req(i_lpddr_ppp_0_pwr_idle_vec_req[0]),
        .i_lpddr_ppp_0_clk(i_lpddr_ppp_0_clk),
        .i_lpddr_ppp_0_clken(i_lpddr_ppp_0_clken),
        .o_lpddr_ppp_0_pwr_idle_val(o_lpddr_ppp_0_pwr_idle_vec_val[1]),
        .o_lpddr_ppp_0_pwr_idle_ack(o_lpddr_ppp_0_pwr_idle_vec_ack[1]),
        .i_lpddr_ppp_0_pwr_idle_req(i_lpddr_ppp_0_pwr_idle_vec_req[1]),
        .i_lpddr_ppp_0_rst_n(i_lpddr_ppp_0_rst_n),
        .o_lpddr_ppp_0_targ_cfg_apb_m_paddr(o_lpddr_ppp_0_targ_cfg_apb_m_paddr),
        .o_lpddr_ppp_0_targ_cfg_apb_m_penable(o_lpddr_ppp_0_targ_cfg_apb_m_penable),
        .o_lpddr_ppp_0_targ_cfg_apb_m_pprot(o_lpddr_ppp_0_targ_cfg_apb_m_pprot),
        .i_lpddr_ppp_0_targ_cfg_apb_m_prdata(i_lpddr_ppp_0_targ_cfg_apb_m_prdata),
        .i_lpddr_ppp_0_targ_cfg_apb_m_pready(i_lpddr_ppp_0_targ_cfg_apb_m_pready),
        .o_lpddr_ppp_0_targ_cfg_apb_m_psel(o_lpddr_ppp_0_targ_cfg_apb_m_psel),
        .i_lpddr_ppp_0_targ_cfg_apb_m_pslverr(i_lpddr_ppp_0_targ_cfg_apb_m_pslverr),
        .o_lpddr_ppp_0_targ_cfg_apb_m_pstrb(o_lpddr_ppp_0_targ_cfg_apb_m_pstrb),
        .o_lpddr_ppp_0_targ_cfg_apb_m_pwdata(o_lpddr_ppp_0_targ_cfg_apb_m_pwdata),
        .o_lpddr_ppp_0_targ_cfg_apb_m_pwrite(o_lpddr_ppp_0_targ_cfg_apb_m_pwrite),
        .o_lpddr_ppp_0_targ_mt_axi_m_araddr(o_lpddr_ppp_0_targ_mt_axi_m_araddr),
        .o_lpddr_ppp_0_targ_mt_axi_m_arburst(o_lpddr_ppp_0_targ_mt_axi_m_arburst),
        .o_lpddr_ppp_0_targ_mt_axi_m_arcache(o_lpddr_ppp_0_targ_mt_axi_m_arcache),
        .o_lpddr_ppp_0_targ_mt_axi_m_arid(o_lpddr_ppp_0_targ_mt_axi_m_arid),
        .o_lpddr_ppp_0_targ_mt_axi_m_arlen(o_lpddr_ppp_0_targ_mt_axi_m_arlen),
        .o_lpddr_ppp_0_targ_mt_axi_m_arlock(o_lpddr_ppp_0_targ_mt_axi_m_arlock),
        .o_lpddr_ppp_0_targ_mt_axi_m_arprot(o_lpddr_ppp_0_targ_mt_axi_m_arprot),
        .o_lpddr_ppp_0_targ_mt_axi_m_arqos(o_lpddr_ppp_0_targ_mt_axi_m_arqos),
        .i_lpddr_ppp_0_targ_mt_axi_m_arready(i_lpddr_ppp_0_targ_mt_axi_m_arready),
        .o_lpddr_ppp_0_targ_mt_axi_m_arsize(o_lpddr_ppp_0_targ_mt_axi_m_arsize),
        .o_lpddr_ppp_0_targ_mt_axi_m_arvalid(o_lpddr_ppp_0_targ_mt_axi_m_arvalid),
        .o_lpddr_ppp_0_targ_mt_axi_m_awaddr(o_lpddr_ppp_0_targ_mt_axi_m_awaddr),
        .o_lpddr_ppp_0_targ_mt_axi_m_awburst(o_lpddr_ppp_0_targ_mt_axi_m_awburst),
        .o_lpddr_ppp_0_targ_mt_axi_m_awcache(o_lpddr_ppp_0_targ_mt_axi_m_awcache),
        .o_lpddr_ppp_0_targ_mt_axi_m_awid(o_lpddr_ppp_0_targ_mt_axi_m_awid),
        .o_lpddr_ppp_0_targ_mt_axi_m_awlen(o_lpddr_ppp_0_targ_mt_axi_m_awlen),
        .o_lpddr_ppp_0_targ_mt_axi_m_awlock(o_lpddr_ppp_0_targ_mt_axi_m_awlock),
        .o_lpddr_ppp_0_targ_mt_axi_m_awprot(o_lpddr_ppp_0_targ_mt_axi_m_awprot),
        .o_lpddr_ppp_0_targ_mt_axi_m_awqos(o_lpddr_ppp_0_targ_mt_axi_m_awqos),
        .i_lpddr_ppp_0_targ_mt_axi_m_awready(i_lpddr_ppp_0_targ_mt_axi_m_awready),
        .o_lpddr_ppp_0_targ_mt_axi_m_awsize(o_lpddr_ppp_0_targ_mt_axi_m_awsize),
        .o_lpddr_ppp_0_targ_mt_axi_m_awvalid(o_lpddr_ppp_0_targ_mt_axi_m_awvalid),
        .i_lpddr_ppp_0_targ_mt_axi_m_bid(i_lpddr_ppp_0_targ_mt_axi_m_bid),
        .o_lpddr_ppp_0_targ_mt_axi_m_bready(o_lpddr_ppp_0_targ_mt_axi_m_bready),
        .i_lpddr_ppp_0_targ_mt_axi_m_bresp(i_lpddr_ppp_0_targ_mt_axi_m_bresp),
        .i_lpddr_ppp_0_targ_mt_axi_m_bvalid(i_lpddr_ppp_0_targ_mt_axi_m_bvalid),
        .i_lpddr_ppp_0_targ_mt_axi_m_rdata(i_lpddr_ppp_0_targ_mt_axi_m_rdata),
        .i_lpddr_ppp_0_targ_mt_axi_m_rid(i_lpddr_ppp_0_targ_mt_axi_m_rid),
        .i_lpddr_ppp_0_targ_mt_axi_m_rlast(i_lpddr_ppp_0_targ_mt_axi_m_rlast),
        .o_lpddr_ppp_0_targ_mt_axi_m_rready(o_lpddr_ppp_0_targ_mt_axi_m_rready),
        .i_lpddr_ppp_0_targ_mt_axi_m_rresp(i_lpddr_ppp_0_targ_mt_axi_m_rresp),
        .i_lpddr_ppp_0_targ_mt_axi_m_rvalid(i_lpddr_ppp_0_targ_mt_axi_m_rvalid),
        .o_lpddr_ppp_0_targ_mt_axi_m_wdata(o_lpddr_ppp_0_targ_mt_axi_m_wdata),
        .o_lpddr_ppp_0_targ_mt_axi_m_wlast(o_lpddr_ppp_0_targ_mt_axi_m_wlast),
        .i_lpddr_ppp_0_targ_mt_axi_m_wready(i_lpddr_ppp_0_targ_mt_axi_m_wready),
        .o_lpddr_ppp_0_targ_mt_axi_m_wstrb(o_lpddr_ppp_0_targ_mt_axi_m_wstrb),
        .o_lpddr_ppp_0_targ_mt_axi_m_wvalid(o_lpddr_ppp_0_targ_mt_axi_m_wvalid),
        .o_lpddr_ppp_0_targ_syscfg_apb_m_paddr(o_lpddr_ppp_0_targ_syscfg_apb_m_paddr),
        .o_lpddr_ppp_0_targ_syscfg_apb_m_penable(o_lpddr_ppp_0_targ_syscfg_apb_m_penable),
        .o_lpddr_ppp_0_targ_syscfg_apb_m_pprot(o_lpddr_ppp_0_targ_syscfg_apb_m_pprot),
        .i_lpddr_ppp_0_targ_syscfg_apb_m_prdata(i_lpddr_ppp_0_targ_syscfg_apb_m_prdata),
        .i_lpddr_ppp_0_targ_syscfg_apb_m_pready(i_lpddr_ppp_0_targ_syscfg_apb_m_pready),
        .o_lpddr_ppp_0_targ_syscfg_apb_m_psel(o_lpddr_ppp_0_targ_syscfg_apb_m_psel),
        .i_lpddr_ppp_0_targ_syscfg_apb_m_pslverr(i_lpddr_ppp_0_targ_syscfg_apb_m_pslverr),
        .o_lpddr_ppp_0_targ_syscfg_apb_m_pstrb(o_lpddr_ppp_0_targ_syscfg_apb_m_pstrb),
        .o_lpddr_ppp_0_targ_syscfg_apb_m_pwdata(o_lpddr_ppp_0_targ_syscfg_apb_m_pwdata),
        .o_lpddr_ppp_0_targ_syscfg_apb_m_pwrite(o_lpddr_ppp_0_targ_syscfg_apb_m_pwrite),
        .i_lpddr_ppp_1_aon_clk(i_lpddr_ppp_1_aon_clk),
        .i_lpddr_ppp_1_aon_rst_n(i_lpddr_ppp_1_aon_rst_n),
        .o_lpddr_ppp_1_cfg_pwr_idle_val(o_lpddr_ppp_1_pwr_idle_vec_val[0]),
        .o_lpddr_ppp_1_cfg_pwr_idle_ack(o_lpddr_ppp_1_pwr_idle_vec_ack[0]),
        .i_lpddr_ppp_1_cfg_pwr_idle_req(i_lpddr_ppp_1_pwr_idle_vec_req[0]),
        .i_lpddr_ppp_1_clk(i_lpddr_ppp_1_clk),
        .i_lpddr_ppp_1_clken(i_lpddr_ppp_1_clken),
        .o_lpddr_ppp_1_pwr_idle_val(o_lpddr_ppp_1_pwr_idle_vec_val[1]),
        .o_lpddr_ppp_1_pwr_idle_ack(o_lpddr_ppp_1_pwr_idle_vec_ack[1]),
        .i_lpddr_ppp_1_pwr_idle_req(i_lpddr_ppp_1_pwr_idle_vec_req[1]),
        .i_lpddr_ppp_1_rst_n(i_lpddr_ppp_1_rst_n),
        .o_lpddr_ppp_1_targ_cfg_apb_m_paddr(o_lpddr_ppp_1_targ_cfg_apb_m_paddr),
        .o_lpddr_ppp_1_targ_cfg_apb_m_penable(o_lpddr_ppp_1_targ_cfg_apb_m_penable),
        .o_lpddr_ppp_1_targ_cfg_apb_m_pprot(o_lpddr_ppp_1_targ_cfg_apb_m_pprot),
        .i_lpddr_ppp_1_targ_cfg_apb_m_prdata(i_lpddr_ppp_1_targ_cfg_apb_m_prdata),
        .i_lpddr_ppp_1_targ_cfg_apb_m_pready(i_lpddr_ppp_1_targ_cfg_apb_m_pready),
        .o_lpddr_ppp_1_targ_cfg_apb_m_psel(o_lpddr_ppp_1_targ_cfg_apb_m_psel),
        .i_lpddr_ppp_1_targ_cfg_apb_m_pslverr(i_lpddr_ppp_1_targ_cfg_apb_m_pslverr),
        .o_lpddr_ppp_1_targ_cfg_apb_m_pstrb(o_lpddr_ppp_1_targ_cfg_apb_m_pstrb),
        .o_lpddr_ppp_1_targ_cfg_apb_m_pwdata(o_lpddr_ppp_1_targ_cfg_apb_m_pwdata),
        .o_lpddr_ppp_1_targ_cfg_apb_m_pwrite(o_lpddr_ppp_1_targ_cfg_apb_m_pwrite),
        .o_lpddr_ppp_1_targ_mt_axi_m_araddr(o_lpddr_ppp_1_targ_mt_axi_m_araddr),
        .o_lpddr_ppp_1_targ_mt_axi_m_arburst(o_lpddr_ppp_1_targ_mt_axi_m_arburst),
        .o_lpddr_ppp_1_targ_mt_axi_m_arcache(o_lpddr_ppp_1_targ_mt_axi_m_arcache),
        .o_lpddr_ppp_1_targ_mt_axi_m_arid(o_lpddr_ppp_1_targ_mt_axi_m_arid),
        .o_lpddr_ppp_1_targ_mt_axi_m_arlen(o_lpddr_ppp_1_targ_mt_axi_m_arlen),
        .o_lpddr_ppp_1_targ_mt_axi_m_arlock(o_lpddr_ppp_1_targ_mt_axi_m_arlock),
        .o_lpddr_ppp_1_targ_mt_axi_m_arprot(o_lpddr_ppp_1_targ_mt_axi_m_arprot),
        .o_lpddr_ppp_1_targ_mt_axi_m_arqos(o_lpddr_ppp_1_targ_mt_axi_m_arqos),
        .i_lpddr_ppp_1_targ_mt_axi_m_arready(i_lpddr_ppp_1_targ_mt_axi_m_arready),
        .o_lpddr_ppp_1_targ_mt_axi_m_arsize(o_lpddr_ppp_1_targ_mt_axi_m_arsize),
        .o_lpddr_ppp_1_targ_mt_axi_m_arvalid(o_lpddr_ppp_1_targ_mt_axi_m_arvalid),
        .o_lpddr_ppp_1_targ_mt_axi_m_awaddr(o_lpddr_ppp_1_targ_mt_axi_m_awaddr),
        .o_lpddr_ppp_1_targ_mt_axi_m_awburst(o_lpddr_ppp_1_targ_mt_axi_m_awburst),
        .o_lpddr_ppp_1_targ_mt_axi_m_awcache(o_lpddr_ppp_1_targ_mt_axi_m_awcache),
        .o_lpddr_ppp_1_targ_mt_axi_m_awid(o_lpddr_ppp_1_targ_mt_axi_m_awid),
        .o_lpddr_ppp_1_targ_mt_axi_m_awlen(o_lpddr_ppp_1_targ_mt_axi_m_awlen),
        .o_lpddr_ppp_1_targ_mt_axi_m_awlock(o_lpddr_ppp_1_targ_mt_axi_m_awlock),
        .o_lpddr_ppp_1_targ_mt_axi_m_awprot(o_lpddr_ppp_1_targ_mt_axi_m_awprot),
        .o_lpddr_ppp_1_targ_mt_axi_m_awqos(o_lpddr_ppp_1_targ_mt_axi_m_awqos),
        .i_lpddr_ppp_1_targ_mt_axi_m_awready(i_lpddr_ppp_1_targ_mt_axi_m_awready),
        .o_lpddr_ppp_1_targ_mt_axi_m_awsize(o_lpddr_ppp_1_targ_mt_axi_m_awsize),
        .o_lpddr_ppp_1_targ_mt_axi_m_awvalid(o_lpddr_ppp_1_targ_mt_axi_m_awvalid),
        .i_lpddr_ppp_1_targ_mt_axi_m_bid(i_lpddr_ppp_1_targ_mt_axi_m_bid),
        .o_lpddr_ppp_1_targ_mt_axi_m_bready(o_lpddr_ppp_1_targ_mt_axi_m_bready),
        .i_lpddr_ppp_1_targ_mt_axi_m_bresp(i_lpddr_ppp_1_targ_mt_axi_m_bresp),
        .i_lpddr_ppp_1_targ_mt_axi_m_bvalid(i_lpddr_ppp_1_targ_mt_axi_m_bvalid),
        .i_lpddr_ppp_1_targ_mt_axi_m_rdata(i_lpddr_ppp_1_targ_mt_axi_m_rdata),
        .i_lpddr_ppp_1_targ_mt_axi_m_rid(i_lpddr_ppp_1_targ_mt_axi_m_rid),
        .i_lpddr_ppp_1_targ_mt_axi_m_rlast(i_lpddr_ppp_1_targ_mt_axi_m_rlast),
        .o_lpddr_ppp_1_targ_mt_axi_m_rready(o_lpddr_ppp_1_targ_mt_axi_m_rready),
        .i_lpddr_ppp_1_targ_mt_axi_m_rresp(i_lpddr_ppp_1_targ_mt_axi_m_rresp),
        .i_lpddr_ppp_1_targ_mt_axi_m_rvalid(i_lpddr_ppp_1_targ_mt_axi_m_rvalid),
        .o_lpddr_ppp_1_targ_mt_axi_m_wdata(o_lpddr_ppp_1_targ_mt_axi_m_wdata),
        .o_lpddr_ppp_1_targ_mt_axi_m_wlast(o_lpddr_ppp_1_targ_mt_axi_m_wlast),
        .i_lpddr_ppp_1_targ_mt_axi_m_wready(i_lpddr_ppp_1_targ_mt_axi_m_wready),
        .o_lpddr_ppp_1_targ_mt_axi_m_wstrb(o_lpddr_ppp_1_targ_mt_axi_m_wstrb),
        .o_lpddr_ppp_1_targ_mt_axi_m_wvalid(o_lpddr_ppp_1_targ_mt_axi_m_wvalid),
        .o_lpddr_ppp_1_targ_syscfg_apb_m_paddr(o_lpddr_ppp_1_targ_syscfg_apb_m_paddr),
        .o_lpddr_ppp_1_targ_syscfg_apb_m_penable(o_lpddr_ppp_1_targ_syscfg_apb_m_penable),
        .o_lpddr_ppp_1_targ_syscfg_apb_m_pprot(o_lpddr_ppp_1_targ_syscfg_apb_m_pprot),
        .i_lpddr_ppp_1_targ_syscfg_apb_m_prdata(i_lpddr_ppp_1_targ_syscfg_apb_m_prdata),
        .i_lpddr_ppp_1_targ_syscfg_apb_m_pready(i_lpddr_ppp_1_targ_syscfg_apb_m_pready),
        .o_lpddr_ppp_1_targ_syscfg_apb_m_psel(o_lpddr_ppp_1_targ_syscfg_apb_m_psel),
        .i_lpddr_ppp_1_targ_syscfg_apb_m_pslverr(i_lpddr_ppp_1_targ_syscfg_apb_m_pslverr),
        .o_lpddr_ppp_1_targ_syscfg_apb_m_pstrb(o_lpddr_ppp_1_targ_syscfg_apb_m_pstrb),
        .o_lpddr_ppp_1_targ_syscfg_apb_m_pwdata(o_lpddr_ppp_1_targ_syscfg_apb_m_pwdata),
        .o_lpddr_ppp_1_targ_syscfg_apb_m_pwrite(o_lpddr_ppp_1_targ_syscfg_apb_m_pwrite),
        .i_lpddr_ppp_2_aon_clk(i_lpddr_ppp_2_aon_clk),
        .i_lpddr_ppp_2_aon_rst_n(i_lpddr_ppp_2_aon_rst_n),
        .o_lpddr_ppp_2_cfg_pwr_idle_val(o_lpddr_ppp_2_pwr_idle_vec_val[0]),
        .o_lpddr_ppp_2_cfg_pwr_idle_ack(o_lpddr_ppp_2_pwr_idle_vec_ack[0]),
        .i_lpddr_ppp_2_cfg_pwr_idle_req(i_lpddr_ppp_2_pwr_idle_vec_req[0]),
        .i_lpddr_ppp_2_clk(i_lpddr_ppp_2_clk),
        .i_lpddr_ppp_2_clken(i_lpddr_ppp_2_clken),
        .o_lpddr_ppp_2_pwr_idle_val(o_lpddr_ppp_2_pwr_idle_vec_val[1]),
        .o_lpddr_ppp_2_pwr_idle_ack(o_lpddr_ppp_2_pwr_idle_vec_ack[1]),
        .i_lpddr_ppp_2_pwr_idle_req(i_lpddr_ppp_2_pwr_idle_vec_req[1]),
        .i_lpddr_ppp_2_rst_n(i_lpddr_ppp_2_rst_n),
        .o_lpddr_ppp_2_targ_cfg_apb_m_paddr(o_lpddr_ppp_2_targ_cfg_apb_m_paddr),
        .o_lpddr_ppp_2_targ_cfg_apb_m_penable(o_lpddr_ppp_2_targ_cfg_apb_m_penable),
        .o_lpddr_ppp_2_targ_cfg_apb_m_pprot(o_lpddr_ppp_2_targ_cfg_apb_m_pprot),
        .i_lpddr_ppp_2_targ_cfg_apb_m_prdata(i_lpddr_ppp_2_targ_cfg_apb_m_prdata),
        .i_lpddr_ppp_2_targ_cfg_apb_m_pready(i_lpddr_ppp_2_targ_cfg_apb_m_pready),
        .o_lpddr_ppp_2_targ_cfg_apb_m_psel(o_lpddr_ppp_2_targ_cfg_apb_m_psel),
        .i_lpddr_ppp_2_targ_cfg_apb_m_pslverr(i_lpddr_ppp_2_targ_cfg_apb_m_pslverr),
        .o_lpddr_ppp_2_targ_cfg_apb_m_pstrb(o_lpddr_ppp_2_targ_cfg_apb_m_pstrb),
        .o_lpddr_ppp_2_targ_cfg_apb_m_pwdata(o_lpddr_ppp_2_targ_cfg_apb_m_pwdata),
        .o_lpddr_ppp_2_targ_cfg_apb_m_pwrite(o_lpddr_ppp_2_targ_cfg_apb_m_pwrite),
        .o_lpddr_ppp_2_targ_mt_axi_m_araddr(o_lpddr_ppp_2_targ_mt_axi_m_araddr),
        .o_lpddr_ppp_2_targ_mt_axi_m_arburst(o_lpddr_ppp_2_targ_mt_axi_m_arburst),
        .o_lpddr_ppp_2_targ_mt_axi_m_arcache(o_lpddr_ppp_2_targ_mt_axi_m_arcache),
        .o_lpddr_ppp_2_targ_mt_axi_m_arid(o_lpddr_ppp_2_targ_mt_axi_m_arid),
        .o_lpddr_ppp_2_targ_mt_axi_m_arlen(o_lpddr_ppp_2_targ_mt_axi_m_arlen),
        .o_lpddr_ppp_2_targ_mt_axi_m_arlock(o_lpddr_ppp_2_targ_mt_axi_m_arlock),
        .o_lpddr_ppp_2_targ_mt_axi_m_arprot(o_lpddr_ppp_2_targ_mt_axi_m_arprot),
        .o_lpddr_ppp_2_targ_mt_axi_m_arqos(o_lpddr_ppp_2_targ_mt_axi_m_arqos),
        .i_lpddr_ppp_2_targ_mt_axi_m_arready(i_lpddr_ppp_2_targ_mt_axi_m_arready),
        .o_lpddr_ppp_2_targ_mt_axi_m_arsize(o_lpddr_ppp_2_targ_mt_axi_m_arsize),
        .o_lpddr_ppp_2_targ_mt_axi_m_arvalid(o_lpddr_ppp_2_targ_mt_axi_m_arvalid),
        .o_lpddr_ppp_2_targ_mt_axi_m_awaddr(o_lpddr_ppp_2_targ_mt_axi_m_awaddr),
        .o_lpddr_ppp_2_targ_mt_axi_m_awburst(o_lpddr_ppp_2_targ_mt_axi_m_awburst),
        .o_lpddr_ppp_2_targ_mt_axi_m_awcache(o_lpddr_ppp_2_targ_mt_axi_m_awcache),
        .o_lpddr_ppp_2_targ_mt_axi_m_awid(o_lpddr_ppp_2_targ_mt_axi_m_awid),
        .o_lpddr_ppp_2_targ_mt_axi_m_awlen(o_lpddr_ppp_2_targ_mt_axi_m_awlen),
        .o_lpddr_ppp_2_targ_mt_axi_m_awlock(o_lpddr_ppp_2_targ_mt_axi_m_awlock),
        .o_lpddr_ppp_2_targ_mt_axi_m_awprot(o_lpddr_ppp_2_targ_mt_axi_m_awprot),
        .o_lpddr_ppp_2_targ_mt_axi_m_awqos(o_lpddr_ppp_2_targ_mt_axi_m_awqos),
        .i_lpddr_ppp_2_targ_mt_axi_m_awready(i_lpddr_ppp_2_targ_mt_axi_m_awready),
        .o_lpddr_ppp_2_targ_mt_axi_m_awsize(o_lpddr_ppp_2_targ_mt_axi_m_awsize),
        .o_lpddr_ppp_2_targ_mt_axi_m_awvalid(o_lpddr_ppp_2_targ_mt_axi_m_awvalid),
        .i_lpddr_ppp_2_targ_mt_axi_m_bid(i_lpddr_ppp_2_targ_mt_axi_m_bid),
        .o_lpddr_ppp_2_targ_mt_axi_m_bready(o_lpddr_ppp_2_targ_mt_axi_m_bready),
        .i_lpddr_ppp_2_targ_mt_axi_m_bresp(i_lpddr_ppp_2_targ_mt_axi_m_bresp),
        .i_lpddr_ppp_2_targ_mt_axi_m_bvalid(i_lpddr_ppp_2_targ_mt_axi_m_bvalid),
        .i_lpddr_ppp_2_targ_mt_axi_m_rdata(i_lpddr_ppp_2_targ_mt_axi_m_rdata),
        .i_lpddr_ppp_2_targ_mt_axi_m_rid(i_lpddr_ppp_2_targ_mt_axi_m_rid),
        .i_lpddr_ppp_2_targ_mt_axi_m_rlast(i_lpddr_ppp_2_targ_mt_axi_m_rlast),
        .o_lpddr_ppp_2_targ_mt_axi_m_rready(o_lpddr_ppp_2_targ_mt_axi_m_rready),
        .i_lpddr_ppp_2_targ_mt_axi_m_rresp(i_lpddr_ppp_2_targ_mt_axi_m_rresp),
        .i_lpddr_ppp_2_targ_mt_axi_m_rvalid(i_lpddr_ppp_2_targ_mt_axi_m_rvalid),
        .o_lpddr_ppp_2_targ_mt_axi_m_wdata(o_lpddr_ppp_2_targ_mt_axi_m_wdata),
        .o_lpddr_ppp_2_targ_mt_axi_m_wlast(o_lpddr_ppp_2_targ_mt_axi_m_wlast),
        .i_lpddr_ppp_2_targ_mt_axi_m_wready(i_lpddr_ppp_2_targ_mt_axi_m_wready),
        .o_lpddr_ppp_2_targ_mt_axi_m_wstrb(o_lpddr_ppp_2_targ_mt_axi_m_wstrb),
        .o_lpddr_ppp_2_targ_mt_axi_m_wvalid(o_lpddr_ppp_2_targ_mt_axi_m_wvalid),
        .o_lpddr_ppp_2_targ_syscfg_apb_m_paddr(o_lpddr_ppp_2_targ_syscfg_apb_m_paddr),
        .o_lpddr_ppp_2_targ_syscfg_apb_m_penable(o_lpddr_ppp_2_targ_syscfg_apb_m_penable),
        .o_lpddr_ppp_2_targ_syscfg_apb_m_pprot(o_lpddr_ppp_2_targ_syscfg_apb_m_pprot),
        .i_lpddr_ppp_2_targ_syscfg_apb_m_prdata(i_lpddr_ppp_2_targ_syscfg_apb_m_prdata),
        .i_lpddr_ppp_2_targ_syscfg_apb_m_pready(i_lpddr_ppp_2_targ_syscfg_apb_m_pready),
        .o_lpddr_ppp_2_targ_syscfg_apb_m_psel(o_lpddr_ppp_2_targ_syscfg_apb_m_psel),
        .i_lpddr_ppp_2_targ_syscfg_apb_m_pslverr(i_lpddr_ppp_2_targ_syscfg_apb_m_pslverr),
        .o_lpddr_ppp_2_targ_syscfg_apb_m_pstrb(o_lpddr_ppp_2_targ_syscfg_apb_m_pstrb),
        .o_lpddr_ppp_2_targ_syscfg_apb_m_pwdata(o_lpddr_ppp_2_targ_syscfg_apb_m_pwdata),
        .o_lpddr_ppp_2_targ_syscfg_apb_m_pwrite(o_lpddr_ppp_2_targ_syscfg_apb_m_pwrite),
        .i_lpddr_ppp_3_aon_clk(i_lpddr_ppp_3_aon_clk),
        .i_lpddr_ppp_3_aon_rst_n(i_lpddr_ppp_3_aon_rst_n),
        .o_lpddr_ppp_3_cfg_pwr_idle_val(o_lpddr_ppp_3_pwr_idle_vec_val[0]),
        .o_lpddr_ppp_3_cfg_pwr_idle_ack(o_lpddr_ppp_3_pwr_idle_vec_ack[0]),
        .i_lpddr_ppp_3_cfg_pwr_idle_req(i_lpddr_ppp_3_pwr_idle_vec_req[0]),
        .i_lpddr_ppp_3_clk(i_lpddr_ppp_3_clk),
        .i_lpddr_ppp_3_clken(i_lpddr_ppp_3_clken),
        .o_lpddr_ppp_3_pwr_idle_val(o_lpddr_ppp_3_pwr_idle_vec_val[1]),
        .o_lpddr_ppp_3_pwr_idle_ack(o_lpddr_ppp_3_pwr_idle_vec_ack[1]),
        .i_lpddr_ppp_3_pwr_idle_req(i_lpddr_ppp_3_pwr_idle_vec_req[1]),
        .i_lpddr_ppp_3_rst_n(i_lpddr_ppp_3_rst_n),
        .o_lpddr_ppp_3_targ_cfg_apb_m_paddr(o_lpddr_ppp_3_targ_cfg_apb_m_paddr),
        .o_lpddr_ppp_3_targ_cfg_apb_m_penable(o_lpddr_ppp_3_targ_cfg_apb_m_penable),
        .o_lpddr_ppp_3_targ_cfg_apb_m_pprot(o_lpddr_ppp_3_targ_cfg_apb_m_pprot),
        .i_lpddr_ppp_3_targ_cfg_apb_m_prdata(i_lpddr_ppp_3_targ_cfg_apb_m_prdata),
        .i_lpddr_ppp_3_targ_cfg_apb_m_pready(i_lpddr_ppp_3_targ_cfg_apb_m_pready),
        .o_lpddr_ppp_3_targ_cfg_apb_m_psel(o_lpddr_ppp_3_targ_cfg_apb_m_psel),
        .i_lpddr_ppp_3_targ_cfg_apb_m_pslverr(i_lpddr_ppp_3_targ_cfg_apb_m_pslverr),
        .o_lpddr_ppp_3_targ_cfg_apb_m_pstrb(o_lpddr_ppp_3_targ_cfg_apb_m_pstrb),
        .o_lpddr_ppp_3_targ_cfg_apb_m_pwdata(o_lpddr_ppp_3_targ_cfg_apb_m_pwdata),
        .o_lpddr_ppp_3_targ_cfg_apb_m_pwrite(o_lpddr_ppp_3_targ_cfg_apb_m_pwrite),
        .o_lpddr_ppp_3_targ_mt_axi_m_araddr(o_lpddr_ppp_3_targ_mt_axi_m_araddr),
        .o_lpddr_ppp_3_targ_mt_axi_m_arburst(o_lpddr_ppp_3_targ_mt_axi_m_arburst),
        .o_lpddr_ppp_3_targ_mt_axi_m_arcache(o_lpddr_ppp_3_targ_mt_axi_m_arcache),
        .o_lpddr_ppp_3_targ_mt_axi_m_arid(o_lpddr_ppp_3_targ_mt_axi_m_arid),
        .o_lpddr_ppp_3_targ_mt_axi_m_arlen(o_lpddr_ppp_3_targ_mt_axi_m_arlen),
        .o_lpddr_ppp_3_targ_mt_axi_m_arlock(o_lpddr_ppp_3_targ_mt_axi_m_arlock),
        .o_lpddr_ppp_3_targ_mt_axi_m_arprot(o_lpddr_ppp_3_targ_mt_axi_m_arprot),
        .o_lpddr_ppp_3_targ_mt_axi_m_arqos(o_lpddr_ppp_3_targ_mt_axi_m_arqos),
        .i_lpddr_ppp_3_targ_mt_axi_m_arready(i_lpddr_ppp_3_targ_mt_axi_m_arready),
        .o_lpddr_ppp_3_targ_mt_axi_m_arsize(o_lpddr_ppp_3_targ_mt_axi_m_arsize),
        .o_lpddr_ppp_3_targ_mt_axi_m_arvalid(o_lpddr_ppp_3_targ_mt_axi_m_arvalid),
        .o_lpddr_ppp_3_targ_mt_axi_m_awaddr(o_lpddr_ppp_3_targ_mt_axi_m_awaddr),
        .o_lpddr_ppp_3_targ_mt_axi_m_awburst(o_lpddr_ppp_3_targ_mt_axi_m_awburst),
        .o_lpddr_ppp_3_targ_mt_axi_m_awcache(o_lpddr_ppp_3_targ_mt_axi_m_awcache),
        .o_lpddr_ppp_3_targ_mt_axi_m_awid(o_lpddr_ppp_3_targ_mt_axi_m_awid),
        .o_lpddr_ppp_3_targ_mt_axi_m_awlen(o_lpddr_ppp_3_targ_mt_axi_m_awlen),
        .o_lpddr_ppp_3_targ_mt_axi_m_awlock(o_lpddr_ppp_3_targ_mt_axi_m_awlock),
        .o_lpddr_ppp_3_targ_mt_axi_m_awprot(o_lpddr_ppp_3_targ_mt_axi_m_awprot),
        .o_lpddr_ppp_3_targ_mt_axi_m_awqos(o_lpddr_ppp_3_targ_mt_axi_m_awqos),
        .i_lpddr_ppp_3_targ_mt_axi_m_awready(i_lpddr_ppp_3_targ_mt_axi_m_awready),
        .o_lpddr_ppp_3_targ_mt_axi_m_awsize(o_lpddr_ppp_3_targ_mt_axi_m_awsize),
        .o_lpddr_ppp_3_targ_mt_axi_m_awvalid(o_lpddr_ppp_3_targ_mt_axi_m_awvalid),
        .i_lpddr_ppp_3_targ_mt_axi_m_bid(i_lpddr_ppp_3_targ_mt_axi_m_bid),
        .o_lpddr_ppp_3_targ_mt_axi_m_bready(o_lpddr_ppp_3_targ_mt_axi_m_bready),
        .i_lpddr_ppp_3_targ_mt_axi_m_bresp(i_lpddr_ppp_3_targ_mt_axi_m_bresp),
        .i_lpddr_ppp_3_targ_mt_axi_m_bvalid(i_lpddr_ppp_3_targ_mt_axi_m_bvalid),
        .i_lpddr_ppp_3_targ_mt_axi_m_rdata(i_lpddr_ppp_3_targ_mt_axi_m_rdata),
        .i_lpddr_ppp_3_targ_mt_axi_m_rid(i_lpddr_ppp_3_targ_mt_axi_m_rid),
        .i_lpddr_ppp_3_targ_mt_axi_m_rlast(i_lpddr_ppp_3_targ_mt_axi_m_rlast),
        .o_lpddr_ppp_3_targ_mt_axi_m_rready(o_lpddr_ppp_3_targ_mt_axi_m_rready),
        .i_lpddr_ppp_3_targ_mt_axi_m_rresp(i_lpddr_ppp_3_targ_mt_axi_m_rresp),
        .i_lpddr_ppp_3_targ_mt_axi_m_rvalid(i_lpddr_ppp_3_targ_mt_axi_m_rvalid),
        .o_lpddr_ppp_3_targ_mt_axi_m_wdata(o_lpddr_ppp_3_targ_mt_axi_m_wdata),
        .o_lpddr_ppp_3_targ_mt_axi_m_wlast(o_lpddr_ppp_3_targ_mt_axi_m_wlast),
        .i_lpddr_ppp_3_targ_mt_axi_m_wready(i_lpddr_ppp_3_targ_mt_axi_m_wready),
        .o_lpddr_ppp_3_targ_mt_axi_m_wstrb(o_lpddr_ppp_3_targ_mt_axi_m_wstrb),
        .o_lpddr_ppp_3_targ_mt_axi_m_wvalid(o_lpddr_ppp_3_targ_mt_axi_m_wvalid),
        .o_lpddr_ppp_3_targ_syscfg_apb_m_paddr(o_lpddr_ppp_3_targ_syscfg_apb_m_paddr),
        .o_lpddr_ppp_3_targ_syscfg_apb_m_penable(o_lpddr_ppp_3_targ_syscfg_apb_m_penable),
        .o_lpddr_ppp_3_targ_syscfg_apb_m_pprot(o_lpddr_ppp_3_targ_syscfg_apb_m_pprot),
        .i_lpddr_ppp_3_targ_syscfg_apb_m_prdata(i_lpddr_ppp_3_targ_syscfg_apb_m_prdata),
        .i_lpddr_ppp_3_targ_syscfg_apb_m_pready(i_lpddr_ppp_3_targ_syscfg_apb_m_pready),
        .o_lpddr_ppp_3_targ_syscfg_apb_m_psel(o_lpddr_ppp_3_targ_syscfg_apb_m_psel),
        .i_lpddr_ppp_3_targ_syscfg_apb_m_pslverr(i_lpddr_ppp_3_targ_syscfg_apb_m_pslverr),
        .o_lpddr_ppp_3_targ_syscfg_apb_m_pstrb(o_lpddr_ppp_3_targ_syscfg_apb_m_pstrb),
        .o_lpddr_ppp_3_targ_syscfg_apb_m_pwdata(o_lpddr_ppp_3_targ_syscfg_apb_m_pwdata),
        .o_lpddr_ppp_3_targ_syscfg_apb_m_pwrite(o_lpddr_ppp_3_targ_syscfg_apb_m_pwrite),
        .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
        .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
        .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
        .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
        .i_noc_clk(i_noc_clk),
        .i_noc_rst_n(i_noc_rst_n),
        .i_soc_periph_aon_clk(i_soc_periph_aon_clk),
        .i_soc_periph_aon_rst_n(i_soc_periph_aon_rst_n),
        .i_soc_periph_clk(i_soc_periph_clk),
        .i_soc_periph_clken(i_soc_periph_clken),
        .i_soc_periph_init_lt_axi_s_araddr(i_soc_periph_init_lt_axi_s_araddr),
        .i_soc_periph_init_lt_axi_s_arburst(i_soc_periph_init_lt_axi_s_arburst),
        .i_soc_periph_init_lt_axi_s_arcache(i_soc_periph_init_lt_axi_s_arcache),
        .i_soc_periph_init_lt_axi_s_arid(i_soc_periph_init_lt_axi_s_arid),
        .i_soc_periph_init_lt_axi_s_arlen(i_soc_periph_init_lt_axi_s_arlen),
        .i_soc_periph_init_lt_axi_s_arlock(i_soc_periph_init_lt_axi_s_arlock),
        .i_soc_periph_init_lt_axi_s_arprot(i_soc_periph_init_lt_axi_s_arprot),
        .i_soc_periph_init_lt_axi_s_arqos(i_soc_periph_init_lt_axi_s_arqos),
        .o_soc_periph_init_lt_axi_s_arready(o_soc_periph_init_lt_axi_s_arready),
        .i_soc_periph_init_lt_axi_s_arsize(i_soc_periph_init_lt_axi_s_arsize),
        .i_soc_periph_init_lt_axi_s_arvalid(i_soc_periph_init_lt_axi_s_arvalid),
        .i_soc_periph_init_lt_axi_s_awaddr(i_soc_periph_init_lt_axi_s_awaddr),
        .i_soc_periph_init_lt_axi_s_awburst(i_soc_periph_init_lt_axi_s_awburst),
        .i_soc_periph_init_lt_axi_s_awcache(i_soc_periph_init_lt_axi_s_awcache),
        .i_soc_periph_init_lt_axi_s_awid(i_soc_periph_init_lt_axi_s_awid),
        .i_soc_periph_init_lt_axi_s_awlen(i_soc_periph_init_lt_axi_s_awlen),
        .i_soc_periph_init_lt_axi_s_awlock(i_soc_periph_init_lt_axi_s_awlock),
        .i_soc_periph_init_lt_axi_s_awprot(i_soc_periph_init_lt_axi_s_awprot),
        .i_soc_periph_init_lt_axi_s_awqos(i_soc_periph_init_lt_axi_s_awqos),
        .o_soc_periph_init_lt_axi_s_awready(o_soc_periph_init_lt_axi_s_awready),
        .i_soc_periph_init_lt_axi_s_awsize(i_soc_periph_init_lt_axi_s_awsize),
        .i_soc_periph_init_lt_axi_s_awvalid(i_soc_periph_init_lt_axi_s_awvalid),
        .o_soc_periph_init_lt_axi_s_bid(o_soc_periph_init_lt_axi_s_bid),
        .i_soc_periph_init_lt_axi_s_bready(i_soc_periph_init_lt_axi_s_bready),
        .o_soc_periph_init_lt_axi_s_bresp(o_soc_periph_init_lt_axi_s_bresp),
        .o_soc_periph_init_lt_axi_s_bvalid(o_soc_periph_init_lt_axi_s_bvalid),
        .o_soc_periph_init_lt_axi_s_rdata(o_soc_periph_init_lt_axi_s_rdata),
        .o_soc_periph_init_lt_axi_s_rid(o_soc_periph_init_lt_axi_s_rid),
        .o_soc_periph_init_lt_axi_s_rlast(o_soc_periph_init_lt_axi_s_rlast),
        .i_soc_periph_init_lt_axi_s_rready(i_soc_periph_init_lt_axi_s_rready),
        .o_soc_periph_init_lt_axi_s_rresp(o_soc_periph_init_lt_axi_s_rresp),
        .o_soc_periph_init_lt_axi_s_rvalid(o_soc_periph_init_lt_axi_s_rvalid),
        .i_soc_periph_init_lt_axi_s_wdata(i_soc_periph_init_lt_axi_s_wdata),
        .i_soc_periph_init_lt_axi_s_wlast(i_soc_periph_init_lt_axi_s_wlast),
        .o_soc_periph_init_lt_axi_s_wready(o_soc_periph_init_lt_axi_s_wready),
        .i_soc_periph_init_lt_axi_s_wstrb(i_soc_periph_init_lt_axi_s_wstrb),
        .i_soc_periph_init_lt_axi_s_wvalid(i_soc_periph_init_lt_axi_s_wvalid),
        .o_soc_periph_pwr_idle_val(o_soc_periph_pwr_idle_val),
        .o_soc_periph_pwr_idle_ack(o_soc_periph_pwr_idle_ack),
        .i_soc_periph_pwr_idle_req(i_soc_periph_pwr_idle_req),
        .i_soc_periph_rst_n(i_soc_periph_rst_n),
        .o_soc_periph_targ_lt_axi_m_araddr(o_soc_periph_targ_lt_axi_m_araddr),
        .o_soc_periph_targ_lt_axi_m_arburst(o_soc_periph_targ_lt_axi_m_arburst),
        .o_soc_periph_targ_lt_axi_m_arcache(o_soc_periph_targ_lt_axi_m_arcache),
        .o_soc_periph_targ_lt_axi_m_arid(o_soc_periph_targ_lt_axi_m_arid),
        .o_soc_periph_targ_lt_axi_m_arlen(o_soc_periph_targ_lt_axi_m_arlen),
        .o_soc_periph_targ_lt_axi_m_arlock(o_soc_periph_targ_lt_axi_m_arlock),
        .o_soc_periph_targ_lt_axi_m_arprot(o_soc_periph_targ_lt_axi_m_arprot),
        .o_soc_periph_targ_lt_axi_m_arqos(o_soc_periph_targ_lt_axi_m_arqos),
        .i_soc_periph_targ_lt_axi_m_arready(i_soc_periph_targ_lt_axi_m_arready),
        .o_soc_periph_targ_lt_axi_m_arsize(o_soc_periph_targ_lt_axi_m_arsize),
        .o_soc_periph_targ_lt_axi_m_arvalid(o_soc_periph_targ_lt_axi_m_arvalid),
        .o_soc_periph_targ_lt_axi_m_awaddr(o_soc_periph_targ_lt_axi_m_awaddr),
        .o_soc_periph_targ_lt_axi_m_awburst(o_soc_periph_targ_lt_axi_m_awburst),
        .o_soc_periph_targ_lt_axi_m_awcache(o_soc_periph_targ_lt_axi_m_awcache),
        .o_soc_periph_targ_lt_axi_m_awid(o_soc_periph_targ_lt_axi_m_awid),
        .o_soc_periph_targ_lt_axi_m_awlen(o_soc_periph_targ_lt_axi_m_awlen),
        .o_soc_periph_targ_lt_axi_m_awlock(o_soc_periph_targ_lt_axi_m_awlock),
        .o_soc_periph_targ_lt_axi_m_awprot(o_soc_periph_targ_lt_axi_m_awprot),
        .o_soc_periph_targ_lt_axi_m_awqos(o_soc_periph_targ_lt_axi_m_awqos),
        .i_soc_periph_targ_lt_axi_m_awready(i_soc_periph_targ_lt_axi_m_awready),
        .o_soc_periph_targ_lt_axi_m_awsize(o_soc_periph_targ_lt_axi_m_awsize),
        .o_soc_periph_targ_lt_axi_m_awvalid(o_soc_periph_targ_lt_axi_m_awvalid),
        .i_soc_periph_targ_lt_axi_m_bid(i_soc_periph_targ_lt_axi_m_bid),
        .o_soc_periph_targ_lt_axi_m_bready(o_soc_periph_targ_lt_axi_m_bready),
        .i_soc_periph_targ_lt_axi_m_bresp(i_soc_periph_targ_lt_axi_m_bresp),
        .i_soc_periph_targ_lt_axi_m_bvalid(i_soc_periph_targ_lt_axi_m_bvalid),
        .i_soc_periph_targ_lt_axi_m_rdata(i_soc_periph_targ_lt_axi_m_rdata),
        .i_soc_periph_targ_lt_axi_m_rid(i_soc_periph_targ_lt_axi_m_rid),
        .i_soc_periph_targ_lt_axi_m_rlast(i_soc_periph_targ_lt_axi_m_rlast),
        .o_soc_periph_targ_lt_axi_m_rready(o_soc_periph_targ_lt_axi_m_rready),
        .i_soc_periph_targ_lt_axi_m_rresp(i_soc_periph_targ_lt_axi_m_rresp),
        .i_soc_periph_targ_lt_axi_m_rvalid(i_soc_periph_targ_lt_axi_m_rvalid),
        .o_soc_periph_targ_lt_axi_m_wdata(o_soc_periph_targ_lt_axi_m_wdata),
        .o_soc_periph_targ_lt_axi_m_wlast(o_soc_periph_targ_lt_axi_m_wlast),
        .i_soc_periph_targ_lt_axi_m_wready(i_soc_periph_targ_lt_axi_m_wready),
        .o_soc_periph_targ_lt_axi_m_wstrb(o_soc_periph_targ_lt_axi_m_wstrb),
        .o_soc_periph_targ_lt_axi_m_wvalid(o_soc_periph_targ_lt_axi_m_wvalid),
        .o_soc_periph_targ_syscfg_apb_m_paddr(o_soc_periph_targ_syscfg_apb_m_paddr),
        .o_soc_periph_targ_syscfg_apb_m_penable(o_soc_periph_targ_syscfg_apb_m_penable),
        .o_soc_periph_targ_syscfg_apb_m_pprot(o_soc_periph_targ_syscfg_apb_m_pprot),
        .i_soc_periph_targ_syscfg_apb_m_prdata(i_soc_periph_targ_syscfg_apb_m_prdata),
        .i_soc_periph_targ_syscfg_apb_m_pready(i_soc_periph_targ_syscfg_apb_m_pready),
        .o_soc_periph_targ_syscfg_apb_m_psel(o_soc_periph_targ_syscfg_apb_m_psel),
        .i_soc_periph_targ_syscfg_apb_m_pslverr(i_soc_periph_targ_syscfg_apb_m_pslverr),
        .o_soc_periph_targ_syscfg_apb_m_pstrb(o_soc_periph_targ_syscfg_apb_m_pstrb),
        .o_soc_periph_targ_syscfg_apb_m_pwdata(o_soc_periph_targ_syscfg_apb_m_pwdata),
        .o_soc_periph_targ_syscfg_apb_m_pwrite(o_soc_periph_targ_syscfg_apb_m_pwrite),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  )
    );

    // Instance of noc_ddr_west_p
    noc_ddr_west_p ddr_west_p (
        .i_ddr_wpll_aon_clk(i_ddr_wpll_aon_clk),
        .i_ddr_wpll_aon_rst_n(i_ddr_wpll_aon_rst_n),
        .o_ddr_wpll_targ_syscfg_apb_m_paddr(o_ddr_wpll_targ_syscfg_apb_m_paddr),
        .o_ddr_wpll_targ_syscfg_apb_m_penable(o_ddr_wpll_targ_syscfg_apb_m_penable),
        .o_ddr_wpll_targ_syscfg_apb_m_pprot(o_ddr_wpll_targ_syscfg_apb_m_pprot),
        .i_ddr_wpll_targ_syscfg_apb_m_prdata(i_ddr_wpll_targ_syscfg_apb_m_prdata),
        .i_ddr_wpll_targ_syscfg_apb_m_pready(i_ddr_wpll_targ_syscfg_apb_m_pready),
        .o_ddr_wpll_targ_syscfg_apb_m_psel(o_ddr_wpll_targ_syscfg_apb_m_psel),
        .i_ddr_wpll_targ_syscfg_apb_m_pslverr(i_ddr_wpll_targ_syscfg_apb_m_pslverr),
        .o_ddr_wpll_targ_syscfg_apb_m_pstrb(o_ddr_wpll_targ_syscfg_apb_m_pstrb),
        .o_ddr_wpll_targ_syscfg_apb_m_pwdata(o_ddr_wpll_targ_syscfg_apb_m_pwdata),
        .o_ddr_wpll_targ_syscfg_apb_m_pwrite(o_ddr_wpll_targ_syscfg_apb_m_pwrite),
        .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data),
        .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head),
        .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy),
        .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail),
        .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld),
        .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data),
        .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head),
        .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy),
        .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail),
        .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld),
        .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data),
        .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head),
        .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy),
        .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail),
        .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld),
        .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data),
        .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head),
        .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy),
        .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail),
        .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld),
        .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data),
        .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head),
        .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy),
        .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail),
        .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld),
        .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data),
        .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head),
        .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy),
        .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail),
        .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld),
        .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data),
        .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head),
        .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy),
        .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail),
        .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld),
        .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data),
        .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head),
        .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy),
        .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail),
        .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld),
        .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data),
        .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head),
        .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy),
        .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail),
        .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld),
        .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data),
        .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head),
        .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy),
        .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail),
        .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld),
        .i_lpddr_graph_0_aon_clk(i_lpddr_graph_0_aon_clk),
        .i_lpddr_graph_0_aon_rst_n(i_lpddr_graph_0_aon_rst_n),
        .o_lpddr_graph_0_cfg_pwr_idle_val(o_lpddr_graph_0_pwr_idle_vec_val[0]),
        .o_lpddr_graph_0_cfg_pwr_idle_ack(o_lpddr_graph_0_pwr_idle_vec_ack[0]),
        .i_lpddr_graph_0_cfg_pwr_idle_req(i_lpddr_graph_0_pwr_idle_vec_req[0]),
        .i_lpddr_graph_0_clk(i_lpddr_graph_0_clk),
        .i_lpddr_graph_0_clken(i_lpddr_graph_0_clken),
        .o_lpddr_graph_0_pwr_idle_val(o_lpddr_graph_0_pwr_idle_vec_val[1]),
        .o_lpddr_graph_0_pwr_idle_ack(o_lpddr_graph_0_pwr_idle_vec_ack[1]),
        .i_lpddr_graph_0_pwr_idle_req(i_lpddr_graph_0_pwr_idle_vec_req[1]),
        .i_lpddr_graph_0_rst_n(i_lpddr_graph_0_rst_n),
        .o_lpddr_graph_0_targ_cfg_apb_m_paddr(o_lpddr_graph_0_targ_cfg_apb_m_paddr),
        .o_lpddr_graph_0_targ_cfg_apb_m_penable(o_lpddr_graph_0_targ_cfg_apb_m_penable),
        .o_lpddr_graph_0_targ_cfg_apb_m_pprot(o_lpddr_graph_0_targ_cfg_apb_m_pprot),
        .i_lpddr_graph_0_targ_cfg_apb_m_prdata(i_lpddr_graph_0_targ_cfg_apb_m_prdata),
        .i_lpddr_graph_0_targ_cfg_apb_m_pready(i_lpddr_graph_0_targ_cfg_apb_m_pready),
        .o_lpddr_graph_0_targ_cfg_apb_m_psel(o_lpddr_graph_0_targ_cfg_apb_m_psel),
        .i_lpddr_graph_0_targ_cfg_apb_m_pslverr(i_lpddr_graph_0_targ_cfg_apb_m_pslverr),
        .o_lpddr_graph_0_targ_cfg_apb_m_pstrb(o_lpddr_graph_0_targ_cfg_apb_m_pstrb),
        .o_lpddr_graph_0_targ_cfg_apb_m_pwdata(o_lpddr_graph_0_targ_cfg_apb_m_pwdata),
        .o_lpddr_graph_0_targ_cfg_apb_m_pwrite(o_lpddr_graph_0_targ_cfg_apb_m_pwrite),
        .o_lpddr_graph_0_targ_ht_axi_m_araddr(o_lpddr_graph_0_targ_ht_axi_m_araddr),
        .o_lpddr_graph_0_targ_ht_axi_m_arburst(o_lpddr_graph_0_targ_ht_axi_m_arburst),
        .o_lpddr_graph_0_targ_ht_axi_m_arcache(o_lpddr_graph_0_targ_ht_axi_m_arcache),
        .o_lpddr_graph_0_targ_ht_axi_m_arid(o_lpddr_graph_0_targ_ht_axi_m_arid),
        .o_lpddr_graph_0_targ_ht_axi_m_arlen(o_lpddr_graph_0_targ_ht_axi_m_arlen),
        .o_lpddr_graph_0_targ_ht_axi_m_arlock(o_lpddr_graph_0_targ_ht_axi_m_arlock),
        .o_lpddr_graph_0_targ_ht_axi_m_arprot(o_lpddr_graph_0_targ_ht_axi_m_arprot),
        .o_lpddr_graph_0_targ_ht_axi_m_arqos(o_lpddr_graph_0_targ_ht_axi_m_arqos),
        .i_lpddr_graph_0_targ_ht_axi_m_arready(i_lpddr_graph_0_targ_ht_axi_m_arready),
        .o_lpddr_graph_0_targ_ht_axi_m_arsize(o_lpddr_graph_0_targ_ht_axi_m_arsize),
        .o_lpddr_graph_0_targ_ht_axi_m_arvalid(o_lpddr_graph_0_targ_ht_axi_m_arvalid),
        .o_lpddr_graph_0_targ_ht_axi_m_awaddr(o_lpddr_graph_0_targ_ht_axi_m_awaddr),
        .o_lpddr_graph_0_targ_ht_axi_m_awburst(o_lpddr_graph_0_targ_ht_axi_m_awburst),
        .o_lpddr_graph_0_targ_ht_axi_m_awcache(o_lpddr_graph_0_targ_ht_axi_m_awcache),
        .o_lpddr_graph_0_targ_ht_axi_m_awid(o_lpddr_graph_0_targ_ht_axi_m_awid),
        .o_lpddr_graph_0_targ_ht_axi_m_awlen(o_lpddr_graph_0_targ_ht_axi_m_awlen),
        .o_lpddr_graph_0_targ_ht_axi_m_awlock(o_lpddr_graph_0_targ_ht_axi_m_awlock),
        .o_lpddr_graph_0_targ_ht_axi_m_awprot(o_lpddr_graph_0_targ_ht_axi_m_awprot),
        .o_lpddr_graph_0_targ_ht_axi_m_awqos(o_lpddr_graph_0_targ_ht_axi_m_awqos),
        .i_lpddr_graph_0_targ_ht_axi_m_awready(i_lpddr_graph_0_targ_ht_axi_m_awready),
        .o_lpddr_graph_0_targ_ht_axi_m_awsize(o_lpddr_graph_0_targ_ht_axi_m_awsize),
        .o_lpddr_graph_0_targ_ht_axi_m_awvalid(o_lpddr_graph_0_targ_ht_axi_m_awvalid),
        .i_lpddr_graph_0_targ_ht_axi_m_bid(i_lpddr_graph_0_targ_ht_axi_m_bid),
        .o_lpddr_graph_0_targ_ht_axi_m_bready(o_lpddr_graph_0_targ_ht_axi_m_bready),
        .i_lpddr_graph_0_targ_ht_axi_m_bresp(i_lpddr_graph_0_targ_ht_axi_m_bresp),
        .i_lpddr_graph_0_targ_ht_axi_m_bvalid(i_lpddr_graph_0_targ_ht_axi_m_bvalid),
        .i_lpddr_graph_0_targ_ht_axi_m_rdata(i_lpddr_graph_0_targ_ht_axi_m_rdata),
        .i_lpddr_graph_0_targ_ht_axi_m_rid(i_lpddr_graph_0_targ_ht_axi_m_rid),
        .i_lpddr_graph_0_targ_ht_axi_m_rlast(i_lpddr_graph_0_targ_ht_axi_m_rlast),
        .o_lpddr_graph_0_targ_ht_axi_m_rready(o_lpddr_graph_0_targ_ht_axi_m_rready),
        .i_lpddr_graph_0_targ_ht_axi_m_rresp(i_lpddr_graph_0_targ_ht_axi_m_rresp),
        .i_lpddr_graph_0_targ_ht_axi_m_rvalid(i_lpddr_graph_0_targ_ht_axi_m_rvalid),
        .o_lpddr_graph_0_targ_ht_axi_m_wdata(o_lpddr_graph_0_targ_ht_axi_m_wdata),
        .o_lpddr_graph_0_targ_ht_axi_m_wlast(o_lpddr_graph_0_targ_ht_axi_m_wlast),
        .i_lpddr_graph_0_targ_ht_axi_m_wready(i_lpddr_graph_0_targ_ht_axi_m_wready),
        .o_lpddr_graph_0_targ_ht_axi_m_wstrb(o_lpddr_graph_0_targ_ht_axi_m_wstrb),
        .o_lpddr_graph_0_targ_ht_axi_m_wvalid(o_lpddr_graph_0_targ_ht_axi_m_wvalid),
        .o_lpddr_graph_0_targ_syscfg_apb_m_paddr(o_lpddr_graph_0_targ_syscfg_apb_m_paddr),
        .o_lpddr_graph_0_targ_syscfg_apb_m_penable(o_lpddr_graph_0_targ_syscfg_apb_m_penable),
        .o_lpddr_graph_0_targ_syscfg_apb_m_pprot(o_lpddr_graph_0_targ_syscfg_apb_m_pprot),
        .i_lpddr_graph_0_targ_syscfg_apb_m_prdata(i_lpddr_graph_0_targ_syscfg_apb_m_prdata),
        .i_lpddr_graph_0_targ_syscfg_apb_m_pready(i_lpddr_graph_0_targ_syscfg_apb_m_pready),
        .o_lpddr_graph_0_targ_syscfg_apb_m_psel(o_lpddr_graph_0_targ_syscfg_apb_m_psel),
        .i_lpddr_graph_0_targ_syscfg_apb_m_pslverr(i_lpddr_graph_0_targ_syscfg_apb_m_pslverr),
        .o_lpddr_graph_0_targ_syscfg_apb_m_pstrb(o_lpddr_graph_0_targ_syscfg_apb_m_pstrb),
        .o_lpddr_graph_0_targ_syscfg_apb_m_pwdata(o_lpddr_graph_0_targ_syscfg_apb_m_pwdata),
        .o_lpddr_graph_0_targ_syscfg_apb_m_pwrite(o_lpddr_graph_0_targ_syscfg_apb_m_pwrite),
        .i_lpddr_graph_1_aon_clk(i_lpddr_graph_1_aon_clk),
        .i_lpddr_graph_1_aon_rst_n(i_lpddr_graph_1_aon_rst_n),
        .o_lpddr_graph_1_cfg_pwr_idle_val(o_lpddr_graph_1_pwr_idle_vec_val[0]),
        .o_lpddr_graph_1_cfg_pwr_idle_ack(o_lpddr_graph_1_pwr_idle_vec_ack[0]),
        .i_lpddr_graph_1_cfg_pwr_idle_req(i_lpddr_graph_1_pwr_idle_vec_req[0]),
        .i_lpddr_graph_1_clk(i_lpddr_graph_1_clk),
        .i_lpddr_graph_1_clken(i_lpddr_graph_1_clken),
        .o_lpddr_graph_1_pwr_idle_val(o_lpddr_graph_1_pwr_idle_vec_val[1]),
        .o_lpddr_graph_1_pwr_idle_ack(o_lpddr_graph_1_pwr_idle_vec_ack[1]),
        .i_lpddr_graph_1_pwr_idle_req(i_lpddr_graph_1_pwr_idle_vec_req[1]),
        .i_lpddr_graph_1_rst_n(i_lpddr_graph_1_rst_n),
        .o_lpddr_graph_1_targ_cfg_apb_m_paddr(o_lpddr_graph_1_targ_cfg_apb_m_paddr),
        .o_lpddr_graph_1_targ_cfg_apb_m_penable(o_lpddr_graph_1_targ_cfg_apb_m_penable),
        .o_lpddr_graph_1_targ_cfg_apb_m_pprot(o_lpddr_graph_1_targ_cfg_apb_m_pprot),
        .i_lpddr_graph_1_targ_cfg_apb_m_prdata(i_lpddr_graph_1_targ_cfg_apb_m_prdata),
        .i_lpddr_graph_1_targ_cfg_apb_m_pready(i_lpddr_graph_1_targ_cfg_apb_m_pready),
        .o_lpddr_graph_1_targ_cfg_apb_m_psel(o_lpddr_graph_1_targ_cfg_apb_m_psel),
        .i_lpddr_graph_1_targ_cfg_apb_m_pslverr(i_lpddr_graph_1_targ_cfg_apb_m_pslverr),
        .o_lpddr_graph_1_targ_cfg_apb_m_pstrb(o_lpddr_graph_1_targ_cfg_apb_m_pstrb),
        .o_lpddr_graph_1_targ_cfg_apb_m_pwdata(o_lpddr_graph_1_targ_cfg_apb_m_pwdata),
        .o_lpddr_graph_1_targ_cfg_apb_m_pwrite(o_lpddr_graph_1_targ_cfg_apb_m_pwrite),
        .o_lpddr_graph_1_targ_ht_axi_m_araddr(o_lpddr_graph_1_targ_ht_axi_m_araddr),
        .o_lpddr_graph_1_targ_ht_axi_m_arburst(o_lpddr_graph_1_targ_ht_axi_m_arburst),
        .o_lpddr_graph_1_targ_ht_axi_m_arcache(o_lpddr_graph_1_targ_ht_axi_m_arcache),
        .o_lpddr_graph_1_targ_ht_axi_m_arid(o_lpddr_graph_1_targ_ht_axi_m_arid),
        .o_lpddr_graph_1_targ_ht_axi_m_arlen(o_lpddr_graph_1_targ_ht_axi_m_arlen),
        .o_lpddr_graph_1_targ_ht_axi_m_arlock(o_lpddr_graph_1_targ_ht_axi_m_arlock),
        .o_lpddr_graph_1_targ_ht_axi_m_arprot(o_lpddr_graph_1_targ_ht_axi_m_arprot),
        .o_lpddr_graph_1_targ_ht_axi_m_arqos(o_lpddr_graph_1_targ_ht_axi_m_arqos),
        .i_lpddr_graph_1_targ_ht_axi_m_arready(i_lpddr_graph_1_targ_ht_axi_m_arready),
        .o_lpddr_graph_1_targ_ht_axi_m_arsize(o_lpddr_graph_1_targ_ht_axi_m_arsize),
        .o_lpddr_graph_1_targ_ht_axi_m_arvalid(o_lpddr_graph_1_targ_ht_axi_m_arvalid),
        .o_lpddr_graph_1_targ_ht_axi_m_awaddr(o_lpddr_graph_1_targ_ht_axi_m_awaddr),
        .o_lpddr_graph_1_targ_ht_axi_m_awburst(o_lpddr_graph_1_targ_ht_axi_m_awburst),
        .o_lpddr_graph_1_targ_ht_axi_m_awcache(o_lpddr_graph_1_targ_ht_axi_m_awcache),
        .o_lpddr_graph_1_targ_ht_axi_m_awid(o_lpddr_graph_1_targ_ht_axi_m_awid),
        .o_lpddr_graph_1_targ_ht_axi_m_awlen(o_lpddr_graph_1_targ_ht_axi_m_awlen),
        .o_lpddr_graph_1_targ_ht_axi_m_awlock(o_lpddr_graph_1_targ_ht_axi_m_awlock),
        .o_lpddr_graph_1_targ_ht_axi_m_awprot(o_lpddr_graph_1_targ_ht_axi_m_awprot),
        .o_lpddr_graph_1_targ_ht_axi_m_awqos(o_lpddr_graph_1_targ_ht_axi_m_awqos),
        .i_lpddr_graph_1_targ_ht_axi_m_awready(i_lpddr_graph_1_targ_ht_axi_m_awready),
        .o_lpddr_graph_1_targ_ht_axi_m_awsize(o_lpddr_graph_1_targ_ht_axi_m_awsize),
        .o_lpddr_graph_1_targ_ht_axi_m_awvalid(o_lpddr_graph_1_targ_ht_axi_m_awvalid),
        .i_lpddr_graph_1_targ_ht_axi_m_bid(i_lpddr_graph_1_targ_ht_axi_m_bid),
        .o_lpddr_graph_1_targ_ht_axi_m_bready(o_lpddr_graph_1_targ_ht_axi_m_bready),
        .i_lpddr_graph_1_targ_ht_axi_m_bresp(i_lpddr_graph_1_targ_ht_axi_m_bresp),
        .i_lpddr_graph_1_targ_ht_axi_m_bvalid(i_lpddr_graph_1_targ_ht_axi_m_bvalid),
        .i_lpddr_graph_1_targ_ht_axi_m_rdata(i_lpddr_graph_1_targ_ht_axi_m_rdata),
        .i_lpddr_graph_1_targ_ht_axi_m_rid(i_lpddr_graph_1_targ_ht_axi_m_rid),
        .i_lpddr_graph_1_targ_ht_axi_m_rlast(i_lpddr_graph_1_targ_ht_axi_m_rlast),
        .o_lpddr_graph_1_targ_ht_axi_m_rready(o_lpddr_graph_1_targ_ht_axi_m_rready),
        .i_lpddr_graph_1_targ_ht_axi_m_rresp(i_lpddr_graph_1_targ_ht_axi_m_rresp),
        .i_lpddr_graph_1_targ_ht_axi_m_rvalid(i_lpddr_graph_1_targ_ht_axi_m_rvalid),
        .o_lpddr_graph_1_targ_ht_axi_m_wdata(o_lpddr_graph_1_targ_ht_axi_m_wdata),
        .o_lpddr_graph_1_targ_ht_axi_m_wlast(o_lpddr_graph_1_targ_ht_axi_m_wlast),
        .i_lpddr_graph_1_targ_ht_axi_m_wready(i_lpddr_graph_1_targ_ht_axi_m_wready),
        .o_lpddr_graph_1_targ_ht_axi_m_wstrb(o_lpddr_graph_1_targ_ht_axi_m_wstrb),
        .o_lpddr_graph_1_targ_ht_axi_m_wvalid(o_lpddr_graph_1_targ_ht_axi_m_wvalid),
        .o_lpddr_graph_1_targ_syscfg_apb_m_paddr(o_lpddr_graph_1_targ_syscfg_apb_m_paddr),
        .o_lpddr_graph_1_targ_syscfg_apb_m_penable(o_lpddr_graph_1_targ_syscfg_apb_m_penable),
        .o_lpddr_graph_1_targ_syscfg_apb_m_pprot(o_lpddr_graph_1_targ_syscfg_apb_m_pprot),
        .i_lpddr_graph_1_targ_syscfg_apb_m_prdata(i_lpddr_graph_1_targ_syscfg_apb_m_prdata),
        .i_lpddr_graph_1_targ_syscfg_apb_m_pready(i_lpddr_graph_1_targ_syscfg_apb_m_pready),
        .o_lpddr_graph_1_targ_syscfg_apb_m_psel(o_lpddr_graph_1_targ_syscfg_apb_m_psel),
        .i_lpddr_graph_1_targ_syscfg_apb_m_pslverr(i_lpddr_graph_1_targ_syscfg_apb_m_pslverr),
        .o_lpddr_graph_1_targ_syscfg_apb_m_pstrb(o_lpddr_graph_1_targ_syscfg_apb_m_pstrb),
        .o_lpddr_graph_1_targ_syscfg_apb_m_pwdata(o_lpddr_graph_1_targ_syscfg_apb_m_pwdata),
        .o_lpddr_graph_1_targ_syscfg_apb_m_pwrite(o_lpddr_graph_1_targ_syscfg_apb_m_pwrite),
        .i_lpddr_graph_2_aon_clk(i_lpddr_graph_2_aon_clk),
        .i_lpddr_graph_2_aon_rst_n(i_lpddr_graph_2_aon_rst_n),
        .o_lpddr_graph_2_cfg_pwr_idle_val(o_lpddr_graph_2_pwr_idle_vec_val[0]),
        .o_lpddr_graph_2_cfg_pwr_idle_ack(o_lpddr_graph_2_pwr_idle_vec_ack[0]),
        .i_lpddr_graph_2_cfg_pwr_idle_req(i_lpddr_graph_2_pwr_idle_vec_req[0]),
        .i_lpddr_graph_2_clk(i_lpddr_graph_2_clk),
        .i_lpddr_graph_2_clken(i_lpddr_graph_2_clken),
        .o_lpddr_graph_2_pwr_idle_val(o_lpddr_graph_2_pwr_idle_vec_val[1]),
        .o_lpddr_graph_2_pwr_idle_ack(o_lpddr_graph_2_pwr_idle_vec_ack[1]),
        .i_lpddr_graph_2_pwr_idle_req(i_lpddr_graph_2_pwr_idle_vec_req[1]),
        .i_lpddr_graph_2_rst_n(i_lpddr_graph_2_rst_n),
        .o_lpddr_graph_2_targ_cfg_apb_m_paddr(o_lpddr_graph_2_targ_cfg_apb_m_paddr),
        .o_lpddr_graph_2_targ_cfg_apb_m_penable(o_lpddr_graph_2_targ_cfg_apb_m_penable),
        .o_lpddr_graph_2_targ_cfg_apb_m_pprot(o_lpddr_graph_2_targ_cfg_apb_m_pprot),
        .i_lpddr_graph_2_targ_cfg_apb_m_prdata(i_lpddr_graph_2_targ_cfg_apb_m_prdata),
        .i_lpddr_graph_2_targ_cfg_apb_m_pready(i_lpddr_graph_2_targ_cfg_apb_m_pready),
        .o_lpddr_graph_2_targ_cfg_apb_m_psel(o_lpddr_graph_2_targ_cfg_apb_m_psel),
        .i_lpddr_graph_2_targ_cfg_apb_m_pslverr(i_lpddr_graph_2_targ_cfg_apb_m_pslverr),
        .o_lpddr_graph_2_targ_cfg_apb_m_pstrb(o_lpddr_graph_2_targ_cfg_apb_m_pstrb),
        .o_lpddr_graph_2_targ_cfg_apb_m_pwdata(o_lpddr_graph_2_targ_cfg_apb_m_pwdata),
        .o_lpddr_graph_2_targ_cfg_apb_m_pwrite(o_lpddr_graph_2_targ_cfg_apb_m_pwrite),
        .o_lpddr_graph_2_targ_ht_axi_m_araddr(o_lpddr_graph_2_targ_ht_axi_m_araddr),
        .o_lpddr_graph_2_targ_ht_axi_m_arburst(o_lpddr_graph_2_targ_ht_axi_m_arburst),
        .o_lpddr_graph_2_targ_ht_axi_m_arcache(o_lpddr_graph_2_targ_ht_axi_m_arcache),
        .o_lpddr_graph_2_targ_ht_axi_m_arid(o_lpddr_graph_2_targ_ht_axi_m_arid),
        .o_lpddr_graph_2_targ_ht_axi_m_arlen(o_lpddr_graph_2_targ_ht_axi_m_arlen),
        .o_lpddr_graph_2_targ_ht_axi_m_arlock(o_lpddr_graph_2_targ_ht_axi_m_arlock),
        .o_lpddr_graph_2_targ_ht_axi_m_arprot(o_lpddr_graph_2_targ_ht_axi_m_arprot),
        .o_lpddr_graph_2_targ_ht_axi_m_arqos(o_lpddr_graph_2_targ_ht_axi_m_arqos),
        .i_lpddr_graph_2_targ_ht_axi_m_arready(i_lpddr_graph_2_targ_ht_axi_m_arready),
        .o_lpddr_graph_2_targ_ht_axi_m_arsize(o_lpddr_graph_2_targ_ht_axi_m_arsize),
        .o_lpddr_graph_2_targ_ht_axi_m_arvalid(o_lpddr_graph_2_targ_ht_axi_m_arvalid),
        .o_lpddr_graph_2_targ_ht_axi_m_awaddr(o_lpddr_graph_2_targ_ht_axi_m_awaddr),
        .o_lpddr_graph_2_targ_ht_axi_m_awburst(o_lpddr_graph_2_targ_ht_axi_m_awburst),
        .o_lpddr_graph_2_targ_ht_axi_m_awcache(o_lpddr_graph_2_targ_ht_axi_m_awcache),
        .o_lpddr_graph_2_targ_ht_axi_m_awid(o_lpddr_graph_2_targ_ht_axi_m_awid),
        .o_lpddr_graph_2_targ_ht_axi_m_awlen(o_lpddr_graph_2_targ_ht_axi_m_awlen),
        .o_lpddr_graph_2_targ_ht_axi_m_awlock(o_lpddr_graph_2_targ_ht_axi_m_awlock),
        .o_lpddr_graph_2_targ_ht_axi_m_awprot(o_lpddr_graph_2_targ_ht_axi_m_awprot),
        .o_lpddr_graph_2_targ_ht_axi_m_awqos(o_lpddr_graph_2_targ_ht_axi_m_awqos),
        .i_lpddr_graph_2_targ_ht_axi_m_awready(i_lpddr_graph_2_targ_ht_axi_m_awready),
        .o_lpddr_graph_2_targ_ht_axi_m_awsize(o_lpddr_graph_2_targ_ht_axi_m_awsize),
        .o_lpddr_graph_2_targ_ht_axi_m_awvalid(o_lpddr_graph_2_targ_ht_axi_m_awvalid),
        .i_lpddr_graph_2_targ_ht_axi_m_bid(i_lpddr_graph_2_targ_ht_axi_m_bid),
        .o_lpddr_graph_2_targ_ht_axi_m_bready(o_lpddr_graph_2_targ_ht_axi_m_bready),
        .i_lpddr_graph_2_targ_ht_axi_m_bresp(i_lpddr_graph_2_targ_ht_axi_m_bresp),
        .i_lpddr_graph_2_targ_ht_axi_m_bvalid(i_lpddr_graph_2_targ_ht_axi_m_bvalid),
        .i_lpddr_graph_2_targ_ht_axi_m_rdata(i_lpddr_graph_2_targ_ht_axi_m_rdata),
        .i_lpddr_graph_2_targ_ht_axi_m_rid(i_lpddr_graph_2_targ_ht_axi_m_rid),
        .i_lpddr_graph_2_targ_ht_axi_m_rlast(i_lpddr_graph_2_targ_ht_axi_m_rlast),
        .o_lpddr_graph_2_targ_ht_axi_m_rready(o_lpddr_graph_2_targ_ht_axi_m_rready),
        .i_lpddr_graph_2_targ_ht_axi_m_rresp(i_lpddr_graph_2_targ_ht_axi_m_rresp),
        .i_lpddr_graph_2_targ_ht_axi_m_rvalid(i_lpddr_graph_2_targ_ht_axi_m_rvalid),
        .o_lpddr_graph_2_targ_ht_axi_m_wdata(o_lpddr_graph_2_targ_ht_axi_m_wdata),
        .o_lpddr_graph_2_targ_ht_axi_m_wlast(o_lpddr_graph_2_targ_ht_axi_m_wlast),
        .i_lpddr_graph_2_targ_ht_axi_m_wready(i_lpddr_graph_2_targ_ht_axi_m_wready),
        .o_lpddr_graph_2_targ_ht_axi_m_wstrb(o_lpddr_graph_2_targ_ht_axi_m_wstrb),
        .o_lpddr_graph_2_targ_ht_axi_m_wvalid(o_lpddr_graph_2_targ_ht_axi_m_wvalid),
        .o_lpddr_graph_2_targ_syscfg_apb_m_paddr(o_lpddr_graph_2_targ_syscfg_apb_m_paddr),
        .o_lpddr_graph_2_targ_syscfg_apb_m_penable(o_lpddr_graph_2_targ_syscfg_apb_m_penable),
        .o_lpddr_graph_2_targ_syscfg_apb_m_pprot(o_lpddr_graph_2_targ_syscfg_apb_m_pprot),
        .i_lpddr_graph_2_targ_syscfg_apb_m_prdata(i_lpddr_graph_2_targ_syscfg_apb_m_prdata),
        .i_lpddr_graph_2_targ_syscfg_apb_m_pready(i_lpddr_graph_2_targ_syscfg_apb_m_pready),
        .o_lpddr_graph_2_targ_syscfg_apb_m_psel(o_lpddr_graph_2_targ_syscfg_apb_m_psel),
        .i_lpddr_graph_2_targ_syscfg_apb_m_pslverr(i_lpddr_graph_2_targ_syscfg_apb_m_pslverr),
        .o_lpddr_graph_2_targ_syscfg_apb_m_pstrb(o_lpddr_graph_2_targ_syscfg_apb_m_pstrb),
        .o_lpddr_graph_2_targ_syscfg_apb_m_pwdata(o_lpddr_graph_2_targ_syscfg_apb_m_pwdata),
        .o_lpddr_graph_2_targ_syscfg_apb_m_pwrite(o_lpddr_graph_2_targ_syscfg_apb_m_pwrite),
        .i_lpddr_graph_3_aon_clk(i_lpddr_graph_3_aon_clk),
        .i_lpddr_graph_3_aon_rst_n(i_lpddr_graph_3_aon_rst_n),
        .o_lpddr_graph_3_cfg_pwr_idle_val(o_lpddr_graph_3_pwr_idle_vec_val[0]),
        .o_lpddr_graph_3_cfg_pwr_idle_ack(o_lpddr_graph_3_pwr_idle_vec_ack[0]),
        .i_lpddr_graph_3_cfg_pwr_idle_req(i_lpddr_graph_3_pwr_idle_vec_req[0]),
        .i_lpddr_graph_3_clk(i_lpddr_graph_3_clk),
        .i_lpddr_graph_3_clken(i_lpddr_graph_3_clken),
        .o_lpddr_graph_3_pwr_idle_val(o_lpddr_graph_3_pwr_idle_vec_val[1]),
        .o_lpddr_graph_3_pwr_idle_ack(o_lpddr_graph_3_pwr_idle_vec_ack[1]),
        .i_lpddr_graph_3_pwr_idle_req(i_lpddr_graph_3_pwr_idle_vec_req[1]),
        .i_lpddr_graph_3_rst_n(i_lpddr_graph_3_rst_n),
        .o_lpddr_graph_3_targ_cfg_apb_m_paddr(o_lpddr_graph_3_targ_cfg_apb_m_paddr),
        .o_lpddr_graph_3_targ_cfg_apb_m_penable(o_lpddr_graph_3_targ_cfg_apb_m_penable),
        .o_lpddr_graph_3_targ_cfg_apb_m_pprot(o_lpddr_graph_3_targ_cfg_apb_m_pprot),
        .i_lpddr_graph_3_targ_cfg_apb_m_prdata(i_lpddr_graph_3_targ_cfg_apb_m_prdata),
        .i_lpddr_graph_3_targ_cfg_apb_m_pready(i_lpddr_graph_3_targ_cfg_apb_m_pready),
        .o_lpddr_graph_3_targ_cfg_apb_m_psel(o_lpddr_graph_3_targ_cfg_apb_m_psel),
        .i_lpddr_graph_3_targ_cfg_apb_m_pslverr(i_lpddr_graph_3_targ_cfg_apb_m_pslverr),
        .o_lpddr_graph_3_targ_cfg_apb_m_pstrb(o_lpddr_graph_3_targ_cfg_apb_m_pstrb),
        .o_lpddr_graph_3_targ_cfg_apb_m_pwdata(o_lpddr_graph_3_targ_cfg_apb_m_pwdata),
        .o_lpddr_graph_3_targ_cfg_apb_m_pwrite(o_lpddr_graph_3_targ_cfg_apb_m_pwrite),
        .o_lpddr_graph_3_targ_ht_axi_m_araddr(o_lpddr_graph_3_targ_ht_axi_m_araddr),
        .o_lpddr_graph_3_targ_ht_axi_m_arburst(o_lpddr_graph_3_targ_ht_axi_m_arburst),
        .o_lpddr_graph_3_targ_ht_axi_m_arcache(o_lpddr_graph_3_targ_ht_axi_m_arcache),
        .o_lpddr_graph_3_targ_ht_axi_m_arid(o_lpddr_graph_3_targ_ht_axi_m_arid),
        .o_lpddr_graph_3_targ_ht_axi_m_arlen(o_lpddr_graph_3_targ_ht_axi_m_arlen),
        .o_lpddr_graph_3_targ_ht_axi_m_arlock(o_lpddr_graph_3_targ_ht_axi_m_arlock),
        .o_lpddr_graph_3_targ_ht_axi_m_arprot(o_lpddr_graph_3_targ_ht_axi_m_arprot),
        .o_lpddr_graph_3_targ_ht_axi_m_arqos(o_lpddr_graph_3_targ_ht_axi_m_arqos),
        .i_lpddr_graph_3_targ_ht_axi_m_arready(i_lpddr_graph_3_targ_ht_axi_m_arready),
        .o_lpddr_graph_3_targ_ht_axi_m_arsize(o_lpddr_graph_3_targ_ht_axi_m_arsize),
        .o_lpddr_graph_3_targ_ht_axi_m_arvalid(o_lpddr_graph_3_targ_ht_axi_m_arvalid),
        .o_lpddr_graph_3_targ_ht_axi_m_awaddr(o_lpddr_graph_3_targ_ht_axi_m_awaddr),
        .o_lpddr_graph_3_targ_ht_axi_m_awburst(o_lpddr_graph_3_targ_ht_axi_m_awburst),
        .o_lpddr_graph_3_targ_ht_axi_m_awcache(o_lpddr_graph_3_targ_ht_axi_m_awcache),
        .o_lpddr_graph_3_targ_ht_axi_m_awid(o_lpddr_graph_3_targ_ht_axi_m_awid),
        .o_lpddr_graph_3_targ_ht_axi_m_awlen(o_lpddr_graph_3_targ_ht_axi_m_awlen),
        .o_lpddr_graph_3_targ_ht_axi_m_awlock(o_lpddr_graph_3_targ_ht_axi_m_awlock),
        .o_lpddr_graph_3_targ_ht_axi_m_awprot(o_lpddr_graph_3_targ_ht_axi_m_awprot),
        .o_lpddr_graph_3_targ_ht_axi_m_awqos(o_lpddr_graph_3_targ_ht_axi_m_awqos),
        .i_lpddr_graph_3_targ_ht_axi_m_awready(i_lpddr_graph_3_targ_ht_axi_m_awready),
        .o_lpddr_graph_3_targ_ht_axi_m_awsize(o_lpddr_graph_3_targ_ht_axi_m_awsize),
        .o_lpddr_graph_3_targ_ht_axi_m_awvalid(o_lpddr_graph_3_targ_ht_axi_m_awvalid),
        .i_lpddr_graph_3_targ_ht_axi_m_bid(i_lpddr_graph_3_targ_ht_axi_m_bid),
        .o_lpddr_graph_3_targ_ht_axi_m_bready(o_lpddr_graph_3_targ_ht_axi_m_bready),
        .i_lpddr_graph_3_targ_ht_axi_m_bresp(i_lpddr_graph_3_targ_ht_axi_m_bresp),
        .i_lpddr_graph_3_targ_ht_axi_m_bvalid(i_lpddr_graph_3_targ_ht_axi_m_bvalid),
        .i_lpddr_graph_3_targ_ht_axi_m_rdata(i_lpddr_graph_3_targ_ht_axi_m_rdata),
        .i_lpddr_graph_3_targ_ht_axi_m_rid(i_lpddr_graph_3_targ_ht_axi_m_rid),
        .i_lpddr_graph_3_targ_ht_axi_m_rlast(i_lpddr_graph_3_targ_ht_axi_m_rlast),
        .o_lpddr_graph_3_targ_ht_axi_m_rready(o_lpddr_graph_3_targ_ht_axi_m_rready),
        .i_lpddr_graph_3_targ_ht_axi_m_rresp(i_lpddr_graph_3_targ_ht_axi_m_rresp),
        .i_lpddr_graph_3_targ_ht_axi_m_rvalid(i_lpddr_graph_3_targ_ht_axi_m_rvalid),
        .o_lpddr_graph_3_targ_ht_axi_m_wdata(o_lpddr_graph_3_targ_ht_axi_m_wdata),
        .o_lpddr_graph_3_targ_ht_axi_m_wlast(o_lpddr_graph_3_targ_ht_axi_m_wlast),
        .i_lpddr_graph_3_targ_ht_axi_m_wready(i_lpddr_graph_3_targ_ht_axi_m_wready),
        .o_lpddr_graph_3_targ_ht_axi_m_wstrb(o_lpddr_graph_3_targ_ht_axi_m_wstrb),
        .o_lpddr_graph_3_targ_ht_axi_m_wvalid(o_lpddr_graph_3_targ_ht_axi_m_wvalid),
        .o_lpddr_graph_3_targ_syscfg_apb_m_paddr(o_lpddr_graph_3_targ_syscfg_apb_m_paddr),
        .o_lpddr_graph_3_targ_syscfg_apb_m_penable(o_lpddr_graph_3_targ_syscfg_apb_m_penable),
        .o_lpddr_graph_3_targ_syscfg_apb_m_pprot(o_lpddr_graph_3_targ_syscfg_apb_m_pprot),
        .i_lpddr_graph_3_targ_syscfg_apb_m_prdata(i_lpddr_graph_3_targ_syscfg_apb_m_prdata),
        .i_lpddr_graph_3_targ_syscfg_apb_m_pready(i_lpddr_graph_3_targ_syscfg_apb_m_pready),
        .o_lpddr_graph_3_targ_syscfg_apb_m_psel(o_lpddr_graph_3_targ_syscfg_apb_m_psel),
        .i_lpddr_graph_3_targ_syscfg_apb_m_pslverr(i_lpddr_graph_3_targ_syscfg_apb_m_pslverr),
        .o_lpddr_graph_3_targ_syscfg_apb_m_pstrb(o_lpddr_graph_3_targ_syscfg_apb_m_pstrb),
        .o_lpddr_graph_3_targ_syscfg_apb_m_pwdata(o_lpddr_graph_3_targ_syscfg_apb_m_pwdata),
        .o_lpddr_graph_3_targ_syscfg_apb_m_pwrite(o_lpddr_graph_3_targ_syscfg_apb_m_pwrite),
        .i_noc_clk(i_noc_clk),
        .i_noc_rst_n(i_noc_rst_n),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  )
    );

    // Instance of noc_h_east_p
    noc_h_east_p h_east_p (
        .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data),
        .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head),
        .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy),
        .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail),
        .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld),
        .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data),
        .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head),
        .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail),
        .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld),
        .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data),
        .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head),
        .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy),
        .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail),
        .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld),
        .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data),
        .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head),
        .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data),
        .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head),
        .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy),
        .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail),
        .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld),
        .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data),
        .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head),
        .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data),
        .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head),
        .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy),
        .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail),
        .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld),
        .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data),
        .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head),
        .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail),
        .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld),
        .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data),
        .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head),
        .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy),
        .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail),
        .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld),
        .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data),
        .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head),
        .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data),
        .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head),
        .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy),
        .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail),
        .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld),
        .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data),
        .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head),
        .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data),
        .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head),
        .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy),
        .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail),
        .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld),
        .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data),
        .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head),
        .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data),
        .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head),
        .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy),
        .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail),
        .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld),
        .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data),
        .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head),
        .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data),
        .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head),
        .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy),
        .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail),
        .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld),
        .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data),
        .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head),
        .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail),
        .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld),
        .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data),
        .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head),
        .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy),
        .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail),
        .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld),
        .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data),
        .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head),
        .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data),
        .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head),
        .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy),
        .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail),
        .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld),
        .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data),
        .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head),
        .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data),
        .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head),
        .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy),
        .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail),
        .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld),
        .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data),
        .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head),
        .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail),
        .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld),

        .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data),
        .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head),
        .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy),
        .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail),
        .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld),
        .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data),
        .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head),
        .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy),
        .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail),
        .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld),
        .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data),
        .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head),
        .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy),
        .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail),
        .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld),
        .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data),
        .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head),
        .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy),
        .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail),
        .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld),
        .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data),
        .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head),
        .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy),
        .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail),
        .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld),
        .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data),
        .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head),
        .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy),
        .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail),
        .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld),
        .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data),
        .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head),
        .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy),
        .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail),
        .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld),
        .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data),
        .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head),
        .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy),
        .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail),
        .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld),

        .i_noc_clk(i_noc_clk),
        .i_noc_rst_n(i_noc_rst_n),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  )
    );

    // Instance of noc_h_north_p

    noc_h_north_p h_north_p (
        .i_aic_4_aon_clk(i_aic_4_aon_clk),
        .i_aic_4_aon_rst_n(i_aic_4_aon_rst_n),
        .i_aic_4_clk(i_aic_4_clk),
        .i_aic_4_clken(i_aic_4_clken),
        .i_aic_4_init_ht_axi_s_araddr(i_aic_4_init_ht_axi_s_araddr),
        .i_aic_4_init_ht_axi_s_arburst(i_aic_4_init_ht_axi_s_arburst),
        .i_aic_4_init_ht_axi_s_arcache(i_aic_4_init_ht_axi_s_arcache),
        .i_aic_4_init_ht_axi_s_arid(i_aic_4_init_ht_axi_s_arid),
        .i_aic_4_init_ht_axi_s_arlen(i_aic_4_init_ht_axi_s_arlen),
        .i_aic_4_init_ht_axi_s_arlock(i_aic_4_init_ht_axi_s_arlock),
        .i_aic_4_init_ht_axi_s_arprot(i_aic_4_init_ht_axi_s_arprot),
        .o_aic_4_init_ht_axi_s_arready(o_aic_4_init_ht_axi_s_arready),
        .i_aic_4_init_ht_axi_s_arsize(i_aic_4_init_ht_axi_s_arsize),
        .i_aic_4_init_ht_axi_s_arvalid(i_aic_4_init_ht_axi_s_arvalid),
        .o_aic_4_init_ht_axi_s_rdata(o_aic_4_init_ht_axi_s_rdata),
        .o_aic_4_init_ht_axi_s_rid(o_aic_4_init_ht_axi_s_rid),
        .o_aic_4_init_ht_axi_s_rlast(o_aic_4_init_ht_axi_s_rlast),
        .i_aic_4_init_ht_axi_s_rready(i_aic_4_init_ht_axi_s_rready),
        .o_aic_4_init_ht_axi_s_rresp(o_aic_4_init_ht_axi_s_rresp),
        .o_aic_4_init_ht_axi_s_rvalid(o_aic_4_init_ht_axi_s_rvalid),
        .i_aic_4_init_ht_axi_s_awaddr(i_aic_4_init_ht_axi_s_awaddr),
        .i_aic_4_init_ht_axi_s_awburst(i_aic_4_init_ht_axi_s_awburst),
        .i_aic_4_init_ht_axi_s_awcache(i_aic_4_init_ht_axi_s_awcache),
        .i_aic_4_init_ht_axi_s_awid(i_aic_4_init_ht_axi_s_awid),
        .i_aic_4_init_ht_axi_s_awlen(i_aic_4_init_ht_axi_s_awlen),
        .i_aic_4_init_ht_axi_s_awlock(i_aic_4_init_ht_axi_s_awlock),
        .i_aic_4_init_ht_axi_s_awprot(i_aic_4_init_ht_axi_s_awprot),
        .o_aic_4_init_ht_axi_s_awready(o_aic_4_init_ht_axi_s_awready),
        .i_aic_4_init_ht_axi_s_awsize(i_aic_4_init_ht_axi_s_awsize),
        .i_aic_4_init_ht_axi_s_awvalid(i_aic_4_init_ht_axi_s_awvalid),
        .o_aic_4_init_ht_axi_s_bid(o_aic_4_init_ht_axi_s_bid),
        .i_aic_4_init_ht_axi_s_bready(i_aic_4_init_ht_axi_s_bready),
        .o_aic_4_init_ht_axi_s_bresp(o_aic_4_init_ht_axi_s_bresp),
        .o_aic_4_init_ht_axi_s_bvalid(o_aic_4_init_ht_axi_s_bvalid),
        .i_aic_4_init_ht_axi_s_wdata(i_aic_4_init_ht_axi_s_wdata),
        .i_aic_4_init_ht_axi_s_wlast(i_aic_4_init_ht_axi_s_wlast),
        .o_aic_4_init_ht_axi_s_wready(o_aic_4_init_ht_axi_s_wready),
        .i_aic_4_init_ht_axi_s_wstrb(i_aic_4_init_ht_axi_s_wstrb),
        .i_aic_4_init_ht_axi_s_wvalid(i_aic_4_init_ht_axi_s_wvalid),
        .i_aic_4_init_lt_axi_s_araddr(i_aic_4_init_lt_axi_s_araddr),
        .i_aic_4_init_lt_axi_s_arburst(i_aic_4_init_lt_axi_s_arburst),
        .i_aic_4_init_lt_axi_s_arcache(i_aic_4_init_lt_axi_s_arcache),
        .i_aic_4_init_lt_axi_s_arid(i_aic_4_init_lt_axi_s_arid),
        .i_aic_4_init_lt_axi_s_arlen(i_aic_4_init_lt_axi_s_arlen),
        .i_aic_4_init_lt_axi_s_arlock(i_aic_4_init_lt_axi_s_arlock),
        .i_aic_4_init_lt_axi_s_arprot(i_aic_4_init_lt_axi_s_arprot),
        .i_aic_4_init_lt_axi_s_arqos(i_aic_4_init_lt_axi_s_arqos),
        .o_aic_4_init_lt_axi_s_arready(o_aic_4_init_lt_axi_s_arready),
        .i_aic_4_init_lt_axi_s_arsize(i_aic_4_init_lt_axi_s_arsize),
        .i_aic_4_init_lt_axi_s_arvalid(i_aic_4_init_lt_axi_s_arvalid),
        .i_aic_4_init_lt_axi_s_awaddr(i_aic_4_init_lt_axi_s_awaddr),
        .i_aic_4_init_lt_axi_s_awburst(i_aic_4_init_lt_axi_s_awburst),
        .i_aic_4_init_lt_axi_s_awcache(i_aic_4_init_lt_axi_s_awcache),
        .i_aic_4_init_lt_axi_s_awid(i_aic_4_init_lt_axi_s_awid),
        .i_aic_4_init_lt_axi_s_awlen(i_aic_4_init_lt_axi_s_awlen),
        .i_aic_4_init_lt_axi_s_awlock(i_aic_4_init_lt_axi_s_awlock),
        .i_aic_4_init_lt_axi_s_awprot(i_aic_4_init_lt_axi_s_awprot),
        .i_aic_4_init_lt_axi_s_awqos(i_aic_4_init_lt_axi_s_awqos),
        .o_aic_4_init_lt_axi_s_awready(o_aic_4_init_lt_axi_s_awready),
        .i_aic_4_init_lt_axi_s_awsize(i_aic_4_init_lt_axi_s_awsize),
        .i_aic_4_init_lt_axi_s_awvalid(i_aic_4_init_lt_axi_s_awvalid),
        .o_aic_4_init_lt_axi_s_bid(o_aic_4_init_lt_axi_s_bid),
        .i_aic_4_init_lt_axi_s_bready(i_aic_4_init_lt_axi_s_bready),
        .o_aic_4_init_lt_axi_s_bresp(o_aic_4_init_lt_axi_s_bresp),
        .o_aic_4_init_lt_axi_s_bvalid(o_aic_4_init_lt_axi_s_bvalid),
        .o_aic_4_init_lt_axi_s_rdata(o_aic_4_init_lt_axi_s_rdata),
        .o_aic_4_init_lt_axi_s_rid(o_aic_4_init_lt_axi_s_rid),
        .o_aic_4_init_lt_axi_s_rlast(o_aic_4_init_lt_axi_s_rlast),
        .i_aic_4_init_lt_axi_s_rready(i_aic_4_init_lt_axi_s_rready),
        .o_aic_4_init_lt_axi_s_rresp(o_aic_4_init_lt_axi_s_rresp),
        .o_aic_4_init_lt_axi_s_rvalid(o_aic_4_init_lt_axi_s_rvalid),
        .i_aic_4_init_lt_axi_s_wdata(i_aic_4_init_lt_axi_s_wdata),
        .i_aic_4_init_lt_axi_s_wlast(i_aic_4_init_lt_axi_s_wlast),
        .o_aic_4_init_lt_axi_s_wready(o_aic_4_init_lt_axi_s_wready),
        .i_aic_4_init_lt_axi_s_wstrb(i_aic_4_init_lt_axi_s_wstrb),
        .i_aic_4_init_lt_axi_s_wvalid(i_aic_4_init_lt_axi_s_wvalid),
        .o_aic_4_pwr_idle_val(o_aic_4_pwr_idle_val),
        .o_aic_4_pwr_idle_ack(o_aic_4_pwr_idle_ack),
        .i_aic_4_pwr_idle_req(i_aic_4_pwr_idle_req),
        .i_aic_4_rst_n(i_aic_4_rst_n),
        .o_aic_4_targ_lt_axi_m_araddr(o_aic_4_targ_lt_axi_m_araddr),
        .o_aic_4_targ_lt_axi_m_arburst(o_aic_4_targ_lt_axi_m_arburst),
        .o_aic_4_targ_lt_axi_m_arcache(o_aic_4_targ_lt_axi_m_arcache),
        .o_aic_4_targ_lt_axi_m_arid(o_aic_4_targ_lt_axi_m_arid),
        .o_aic_4_targ_lt_axi_m_arlen(o_aic_4_targ_lt_axi_m_arlen),
        .o_aic_4_targ_lt_axi_m_arlock(o_aic_4_targ_lt_axi_m_arlock),
        .o_aic_4_targ_lt_axi_m_arprot(o_aic_4_targ_lt_axi_m_arprot),
        .o_aic_4_targ_lt_axi_m_arqos(o_aic_4_targ_lt_axi_m_arqos),
        .i_aic_4_targ_lt_axi_m_arready(i_aic_4_targ_lt_axi_m_arready),
        .o_aic_4_targ_lt_axi_m_arsize(o_aic_4_targ_lt_axi_m_arsize),
        .o_aic_4_targ_lt_axi_m_arvalid(o_aic_4_targ_lt_axi_m_arvalid),
        .o_aic_4_targ_lt_axi_m_awaddr(o_aic_4_targ_lt_axi_m_awaddr),
        .o_aic_4_targ_lt_axi_m_awburst(o_aic_4_targ_lt_axi_m_awburst),
        .o_aic_4_targ_lt_axi_m_awcache(o_aic_4_targ_lt_axi_m_awcache),
        .o_aic_4_targ_lt_axi_m_awid(o_aic_4_targ_lt_axi_m_awid),
        .o_aic_4_targ_lt_axi_m_awlen(o_aic_4_targ_lt_axi_m_awlen),
        .o_aic_4_targ_lt_axi_m_awlock(o_aic_4_targ_lt_axi_m_awlock),
        .o_aic_4_targ_lt_axi_m_awprot(o_aic_4_targ_lt_axi_m_awprot),
        .o_aic_4_targ_lt_axi_m_awqos(o_aic_4_targ_lt_axi_m_awqos),
        .i_aic_4_targ_lt_axi_m_awready(i_aic_4_targ_lt_axi_m_awready),
        .o_aic_4_targ_lt_axi_m_awsize(o_aic_4_targ_lt_axi_m_awsize),
        .o_aic_4_targ_lt_axi_m_awvalid(o_aic_4_targ_lt_axi_m_awvalid),
        .i_aic_4_targ_lt_axi_m_bid(i_aic_4_targ_lt_axi_m_bid),
        .o_aic_4_targ_lt_axi_m_bready(o_aic_4_targ_lt_axi_m_bready),
        .i_aic_4_targ_lt_axi_m_bresp(i_aic_4_targ_lt_axi_m_bresp),
        .i_aic_4_targ_lt_axi_m_bvalid(i_aic_4_targ_lt_axi_m_bvalid),
        .i_aic_4_targ_lt_axi_m_rdata(i_aic_4_targ_lt_axi_m_rdata),
        .i_aic_4_targ_lt_axi_m_rid(i_aic_4_targ_lt_axi_m_rid),
        .i_aic_4_targ_lt_axi_m_rlast(i_aic_4_targ_lt_axi_m_rlast),
        .o_aic_4_targ_lt_axi_m_rready(o_aic_4_targ_lt_axi_m_rready),
        .i_aic_4_targ_lt_axi_m_rresp(i_aic_4_targ_lt_axi_m_rresp),
        .i_aic_4_targ_lt_axi_m_rvalid(i_aic_4_targ_lt_axi_m_rvalid),
        .o_aic_4_targ_lt_axi_m_wdata(o_aic_4_targ_lt_axi_m_wdata),
        .o_aic_4_targ_lt_axi_m_wlast(o_aic_4_targ_lt_axi_m_wlast),
        .i_aic_4_targ_lt_axi_m_wready(i_aic_4_targ_lt_axi_m_wready),
        .o_aic_4_targ_lt_axi_m_wstrb(o_aic_4_targ_lt_axi_m_wstrb),
        .o_aic_4_targ_lt_axi_m_wvalid(o_aic_4_targ_lt_axi_m_wvalid),
        .o_aic_4_targ_syscfg_apb_m_paddr(o_aic_4_targ_syscfg_apb_m_paddr),
        .o_aic_4_targ_syscfg_apb_m_penable(o_aic_4_targ_syscfg_apb_m_penable),
        .o_aic_4_targ_syscfg_apb_m_pprot(o_aic_4_targ_syscfg_apb_m_pprot),
        .i_aic_4_targ_syscfg_apb_m_prdata(i_aic_4_targ_syscfg_apb_m_prdata),
        .i_aic_4_targ_syscfg_apb_m_pready(i_aic_4_targ_syscfg_apb_m_pready),
        .o_aic_4_targ_syscfg_apb_m_psel(o_aic_4_targ_syscfg_apb_m_psel),
        .i_aic_4_targ_syscfg_apb_m_pslverr(i_aic_4_targ_syscfg_apb_m_pslverr),
        .o_aic_4_targ_syscfg_apb_m_pstrb(o_aic_4_targ_syscfg_apb_m_pstrb),
        .o_aic_4_targ_syscfg_apb_m_pwdata(o_aic_4_targ_syscfg_apb_m_pwdata),
        .o_aic_4_targ_syscfg_apb_m_pwrite(o_aic_4_targ_syscfg_apb_m_pwrite),
        .i_aic_5_aon_clk(i_aic_5_aon_clk),
        .i_aic_5_aon_rst_n(i_aic_5_aon_rst_n),
        .i_aic_5_clk(i_aic_5_clk),
        .i_aic_5_clken(i_aic_5_clken),
        .i_aic_5_init_ht_axi_s_araddr(i_aic_5_init_ht_axi_s_araddr),
        .i_aic_5_init_ht_axi_s_arburst(i_aic_5_init_ht_axi_s_arburst),
        .i_aic_5_init_ht_axi_s_arcache(i_aic_5_init_ht_axi_s_arcache),
        .i_aic_5_init_ht_axi_s_arid(i_aic_5_init_ht_axi_s_arid),
        .i_aic_5_init_ht_axi_s_arlen(i_aic_5_init_ht_axi_s_arlen),
        .i_aic_5_init_ht_axi_s_arlock(i_aic_5_init_ht_axi_s_arlock),
        .i_aic_5_init_ht_axi_s_arprot(i_aic_5_init_ht_axi_s_arprot),
        .o_aic_5_init_ht_axi_s_arready(o_aic_5_init_ht_axi_s_arready),
        .i_aic_5_init_ht_axi_s_arsize(i_aic_5_init_ht_axi_s_arsize),
        .i_aic_5_init_ht_axi_s_arvalid(i_aic_5_init_ht_axi_s_arvalid),
        .o_aic_5_init_ht_axi_s_rdata(o_aic_5_init_ht_axi_s_rdata),
        .o_aic_5_init_ht_axi_s_rid(o_aic_5_init_ht_axi_s_rid),
        .o_aic_5_init_ht_axi_s_rlast(o_aic_5_init_ht_axi_s_rlast),
        .i_aic_5_init_ht_axi_s_rready(i_aic_5_init_ht_axi_s_rready),
        .o_aic_5_init_ht_axi_s_rresp(o_aic_5_init_ht_axi_s_rresp),
        .o_aic_5_init_ht_axi_s_rvalid(o_aic_5_init_ht_axi_s_rvalid),
        .i_aic_5_init_ht_axi_s_awaddr(i_aic_5_init_ht_axi_s_awaddr),
        .i_aic_5_init_ht_axi_s_awburst(i_aic_5_init_ht_axi_s_awburst),
        .i_aic_5_init_ht_axi_s_awcache(i_aic_5_init_ht_axi_s_awcache),
        .i_aic_5_init_ht_axi_s_awid(i_aic_5_init_ht_axi_s_awid),
        .i_aic_5_init_ht_axi_s_awlen(i_aic_5_init_ht_axi_s_awlen),
        .i_aic_5_init_ht_axi_s_awlock(i_aic_5_init_ht_axi_s_awlock),
        .i_aic_5_init_ht_axi_s_awprot(i_aic_5_init_ht_axi_s_awprot),
        .o_aic_5_init_ht_axi_s_awready(o_aic_5_init_ht_axi_s_awready),
        .i_aic_5_init_ht_axi_s_awsize(i_aic_5_init_ht_axi_s_awsize),
        .i_aic_5_init_ht_axi_s_awvalid(i_aic_5_init_ht_axi_s_awvalid),
        .o_aic_5_init_ht_axi_s_bid(o_aic_5_init_ht_axi_s_bid),
        .i_aic_5_init_ht_axi_s_bready(i_aic_5_init_ht_axi_s_bready),
        .o_aic_5_init_ht_axi_s_bresp(o_aic_5_init_ht_axi_s_bresp),
        .o_aic_5_init_ht_axi_s_bvalid(o_aic_5_init_ht_axi_s_bvalid),
        .i_aic_5_init_ht_axi_s_wdata(i_aic_5_init_ht_axi_s_wdata),
        .i_aic_5_init_ht_axi_s_wlast(i_aic_5_init_ht_axi_s_wlast),
        .o_aic_5_init_ht_axi_s_wready(o_aic_5_init_ht_axi_s_wready),
        .i_aic_5_init_ht_axi_s_wstrb(i_aic_5_init_ht_axi_s_wstrb),
        .i_aic_5_init_ht_axi_s_wvalid(i_aic_5_init_ht_axi_s_wvalid),
        .i_aic_5_init_lt_axi_s_araddr(i_aic_5_init_lt_axi_s_araddr),
        .i_aic_5_init_lt_axi_s_arburst(i_aic_5_init_lt_axi_s_arburst),
        .i_aic_5_init_lt_axi_s_arcache(i_aic_5_init_lt_axi_s_arcache),
        .i_aic_5_init_lt_axi_s_arid(i_aic_5_init_lt_axi_s_arid),
        .i_aic_5_init_lt_axi_s_arlen(i_aic_5_init_lt_axi_s_arlen),
        .i_aic_5_init_lt_axi_s_arlock(i_aic_5_init_lt_axi_s_arlock),
        .i_aic_5_init_lt_axi_s_arprot(i_aic_5_init_lt_axi_s_arprot),
        .i_aic_5_init_lt_axi_s_arqos(i_aic_5_init_lt_axi_s_arqos),
        .o_aic_5_init_lt_axi_s_arready(o_aic_5_init_lt_axi_s_arready),
        .i_aic_5_init_lt_axi_s_arsize(i_aic_5_init_lt_axi_s_arsize),
        .i_aic_5_init_lt_axi_s_arvalid(i_aic_5_init_lt_axi_s_arvalid),
        .i_aic_5_init_lt_axi_s_awaddr(i_aic_5_init_lt_axi_s_awaddr),
        .i_aic_5_init_lt_axi_s_awburst(i_aic_5_init_lt_axi_s_awburst),
        .i_aic_5_init_lt_axi_s_awcache(i_aic_5_init_lt_axi_s_awcache),
        .i_aic_5_init_lt_axi_s_awid(i_aic_5_init_lt_axi_s_awid),
        .i_aic_5_init_lt_axi_s_awlen(i_aic_5_init_lt_axi_s_awlen),
        .i_aic_5_init_lt_axi_s_awlock(i_aic_5_init_lt_axi_s_awlock),
        .i_aic_5_init_lt_axi_s_awprot(i_aic_5_init_lt_axi_s_awprot),
        .i_aic_5_init_lt_axi_s_awqos(i_aic_5_init_lt_axi_s_awqos),
        .o_aic_5_init_lt_axi_s_awready(o_aic_5_init_lt_axi_s_awready),
        .i_aic_5_init_lt_axi_s_awsize(i_aic_5_init_lt_axi_s_awsize),
        .i_aic_5_init_lt_axi_s_awvalid(i_aic_5_init_lt_axi_s_awvalid),
        .o_aic_5_init_lt_axi_s_bid(o_aic_5_init_lt_axi_s_bid),
        .i_aic_5_init_lt_axi_s_bready(i_aic_5_init_lt_axi_s_bready),
        .o_aic_5_init_lt_axi_s_bresp(o_aic_5_init_lt_axi_s_bresp),
        .o_aic_5_init_lt_axi_s_bvalid(o_aic_5_init_lt_axi_s_bvalid),
        .o_aic_5_init_lt_axi_s_rdata(o_aic_5_init_lt_axi_s_rdata),
        .o_aic_5_init_lt_axi_s_rid(o_aic_5_init_lt_axi_s_rid),
        .o_aic_5_init_lt_axi_s_rlast(o_aic_5_init_lt_axi_s_rlast),
        .i_aic_5_init_lt_axi_s_rready(i_aic_5_init_lt_axi_s_rready),
        .o_aic_5_init_lt_axi_s_rresp(o_aic_5_init_lt_axi_s_rresp),
        .o_aic_5_init_lt_axi_s_rvalid(o_aic_5_init_lt_axi_s_rvalid),
        .i_aic_5_init_lt_axi_s_wdata(i_aic_5_init_lt_axi_s_wdata),
        .i_aic_5_init_lt_axi_s_wlast(i_aic_5_init_lt_axi_s_wlast),
        .o_aic_5_init_lt_axi_s_wready(o_aic_5_init_lt_axi_s_wready),
        .i_aic_5_init_lt_axi_s_wstrb(i_aic_5_init_lt_axi_s_wstrb),
        .i_aic_5_init_lt_axi_s_wvalid(i_aic_5_init_lt_axi_s_wvalid),
        .o_aic_5_pwr_idle_val(o_aic_5_pwr_idle_val),
        .o_aic_5_pwr_idle_ack(o_aic_5_pwr_idle_ack),
        .i_aic_5_pwr_idle_req(i_aic_5_pwr_idle_req),
        .i_aic_5_rst_n(i_aic_5_rst_n),
        .o_aic_5_targ_lt_axi_m_araddr(o_aic_5_targ_lt_axi_m_araddr),
        .o_aic_5_targ_lt_axi_m_arburst(o_aic_5_targ_lt_axi_m_arburst),
        .o_aic_5_targ_lt_axi_m_arcache(o_aic_5_targ_lt_axi_m_arcache),
        .o_aic_5_targ_lt_axi_m_arid(o_aic_5_targ_lt_axi_m_arid),
        .o_aic_5_targ_lt_axi_m_arlen(o_aic_5_targ_lt_axi_m_arlen),
        .o_aic_5_targ_lt_axi_m_arlock(o_aic_5_targ_lt_axi_m_arlock),
        .o_aic_5_targ_lt_axi_m_arprot(o_aic_5_targ_lt_axi_m_arprot),
        .o_aic_5_targ_lt_axi_m_arqos(o_aic_5_targ_lt_axi_m_arqos),
        .i_aic_5_targ_lt_axi_m_arready(i_aic_5_targ_lt_axi_m_arready),
        .o_aic_5_targ_lt_axi_m_arsize(o_aic_5_targ_lt_axi_m_arsize),
        .o_aic_5_targ_lt_axi_m_arvalid(o_aic_5_targ_lt_axi_m_arvalid),
        .o_aic_5_targ_lt_axi_m_awaddr(o_aic_5_targ_lt_axi_m_awaddr),
        .o_aic_5_targ_lt_axi_m_awburst(o_aic_5_targ_lt_axi_m_awburst),
        .o_aic_5_targ_lt_axi_m_awcache(o_aic_5_targ_lt_axi_m_awcache),
        .o_aic_5_targ_lt_axi_m_awid(o_aic_5_targ_lt_axi_m_awid),
        .o_aic_5_targ_lt_axi_m_awlen(o_aic_5_targ_lt_axi_m_awlen),
        .o_aic_5_targ_lt_axi_m_awlock(o_aic_5_targ_lt_axi_m_awlock),
        .o_aic_5_targ_lt_axi_m_awprot(o_aic_5_targ_lt_axi_m_awprot),
        .o_aic_5_targ_lt_axi_m_awqos(o_aic_5_targ_lt_axi_m_awqos),
        .i_aic_5_targ_lt_axi_m_awready(i_aic_5_targ_lt_axi_m_awready),
        .o_aic_5_targ_lt_axi_m_awsize(o_aic_5_targ_lt_axi_m_awsize),
        .o_aic_5_targ_lt_axi_m_awvalid(o_aic_5_targ_lt_axi_m_awvalid),
        .i_aic_5_targ_lt_axi_m_bid(i_aic_5_targ_lt_axi_m_bid),
        .o_aic_5_targ_lt_axi_m_bready(o_aic_5_targ_lt_axi_m_bready),
        .i_aic_5_targ_lt_axi_m_bresp(i_aic_5_targ_lt_axi_m_bresp),
        .i_aic_5_targ_lt_axi_m_bvalid(i_aic_5_targ_lt_axi_m_bvalid),
        .i_aic_5_targ_lt_axi_m_rdata(i_aic_5_targ_lt_axi_m_rdata),
        .i_aic_5_targ_lt_axi_m_rid(i_aic_5_targ_lt_axi_m_rid),
        .i_aic_5_targ_lt_axi_m_rlast(i_aic_5_targ_lt_axi_m_rlast),
        .o_aic_5_targ_lt_axi_m_rready(o_aic_5_targ_lt_axi_m_rready),
        .i_aic_5_targ_lt_axi_m_rresp(i_aic_5_targ_lt_axi_m_rresp),
        .i_aic_5_targ_lt_axi_m_rvalid(i_aic_5_targ_lt_axi_m_rvalid),
        .o_aic_5_targ_lt_axi_m_wdata(o_aic_5_targ_lt_axi_m_wdata),
        .o_aic_5_targ_lt_axi_m_wlast(o_aic_5_targ_lt_axi_m_wlast),
        .i_aic_5_targ_lt_axi_m_wready(i_aic_5_targ_lt_axi_m_wready),
        .o_aic_5_targ_lt_axi_m_wstrb(o_aic_5_targ_lt_axi_m_wstrb),
        .o_aic_5_targ_lt_axi_m_wvalid(o_aic_5_targ_lt_axi_m_wvalid),
        .o_aic_5_targ_syscfg_apb_m_paddr(o_aic_5_targ_syscfg_apb_m_paddr),
        .o_aic_5_targ_syscfg_apb_m_penable(o_aic_5_targ_syscfg_apb_m_penable),
        .o_aic_5_targ_syscfg_apb_m_pprot(o_aic_5_targ_syscfg_apb_m_pprot),
        .i_aic_5_targ_syscfg_apb_m_prdata(i_aic_5_targ_syscfg_apb_m_prdata),
        .i_aic_5_targ_syscfg_apb_m_pready(i_aic_5_targ_syscfg_apb_m_pready),
        .o_aic_5_targ_syscfg_apb_m_psel(o_aic_5_targ_syscfg_apb_m_psel),
        .i_aic_5_targ_syscfg_apb_m_pslverr(i_aic_5_targ_syscfg_apb_m_pslverr),
        .o_aic_5_targ_syscfg_apb_m_pstrb(o_aic_5_targ_syscfg_apb_m_pstrb),
        .o_aic_5_targ_syscfg_apb_m_pwdata(o_aic_5_targ_syscfg_apb_m_pwdata),
        .o_aic_5_targ_syscfg_apb_m_pwrite(o_aic_5_targ_syscfg_apb_m_pwrite),
        .i_aic_6_aon_clk(i_aic_6_aon_clk),
        .i_aic_6_aon_rst_n(i_aic_6_aon_rst_n),
        .i_aic_6_clk(i_aic_6_clk),
        .i_aic_6_clken(i_aic_6_clken),
        .i_aic_6_init_ht_axi_s_araddr(i_aic_6_init_ht_axi_s_araddr),
        .i_aic_6_init_ht_axi_s_arburst(i_aic_6_init_ht_axi_s_arburst),
        .i_aic_6_init_ht_axi_s_arcache(i_aic_6_init_ht_axi_s_arcache),
        .i_aic_6_init_ht_axi_s_arid(i_aic_6_init_ht_axi_s_arid),
        .i_aic_6_init_ht_axi_s_arlen(i_aic_6_init_ht_axi_s_arlen),
        .i_aic_6_init_ht_axi_s_arlock(i_aic_6_init_ht_axi_s_arlock),
        .i_aic_6_init_ht_axi_s_arprot(i_aic_6_init_ht_axi_s_arprot),
        .o_aic_6_init_ht_axi_s_arready(o_aic_6_init_ht_axi_s_arready),
        .i_aic_6_init_ht_axi_s_arsize(i_aic_6_init_ht_axi_s_arsize),
        .i_aic_6_init_ht_axi_s_arvalid(i_aic_6_init_ht_axi_s_arvalid),
        .o_aic_6_init_ht_axi_s_rdata(o_aic_6_init_ht_axi_s_rdata),
        .o_aic_6_init_ht_axi_s_rid(o_aic_6_init_ht_axi_s_rid),
        .o_aic_6_init_ht_axi_s_rlast(o_aic_6_init_ht_axi_s_rlast),
        .i_aic_6_init_ht_axi_s_rready(i_aic_6_init_ht_axi_s_rready),
        .o_aic_6_init_ht_axi_s_rresp(o_aic_6_init_ht_axi_s_rresp),
        .o_aic_6_init_ht_axi_s_rvalid(o_aic_6_init_ht_axi_s_rvalid),
        .i_aic_6_init_ht_axi_s_awaddr(i_aic_6_init_ht_axi_s_awaddr),
        .i_aic_6_init_ht_axi_s_awburst(i_aic_6_init_ht_axi_s_awburst),
        .i_aic_6_init_ht_axi_s_awcache(i_aic_6_init_ht_axi_s_awcache),
        .i_aic_6_init_ht_axi_s_awid(i_aic_6_init_ht_axi_s_awid),
        .i_aic_6_init_ht_axi_s_awlen(i_aic_6_init_ht_axi_s_awlen),
        .i_aic_6_init_ht_axi_s_awlock(i_aic_6_init_ht_axi_s_awlock),
        .i_aic_6_init_ht_axi_s_awprot(i_aic_6_init_ht_axi_s_awprot),
        .o_aic_6_init_ht_axi_s_awready(o_aic_6_init_ht_axi_s_awready),
        .i_aic_6_init_ht_axi_s_awsize(i_aic_6_init_ht_axi_s_awsize),
        .i_aic_6_init_ht_axi_s_awvalid(i_aic_6_init_ht_axi_s_awvalid),
        .o_aic_6_init_ht_axi_s_bid(o_aic_6_init_ht_axi_s_bid),
        .i_aic_6_init_ht_axi_s_bready(i_aic_6_init_ht_axi_s_bready),
        .o_aic_6_init_ht_axi_s_bresp(o_aic_6_init_ht_axi_s_bresp),
        .o_aic_6_init_ht_axi_s_bvalid(o_aic_6_init_ht_axi_s_bvalid),
        .i_aic_6_init_ht_axi_s_wdata(i_aic_6_init_ht_axi_s_wdata),
        .i_aic_6_init_ht_axi_s_wlast(i_aic_6_init_ht_axi_s_wlast),
        .o_aic_6_init_ht_axi_s_wready(o_aic_6_init_ht_axi_s_wready),
        .i_aic_6_init_ht_axi_s_wstrb(i_aic_6_init_ht_axi_s_wstrb),
        .i_aic_6_init_ht_axi_s_wvalid(i_aic_6_init_ht_axi_s_wvalid),
        .i_aic_6_init_lt_axi_s_araddr(i_aic_6_init_lt_axi_s_araddr),
        .i_aic_6_init_lt_axi_s_arburst(i_aic_6_init_lt_axi_s_arburst),
        .i_aic_6_init_lt_axi_s_arcache(i_aic_6_init_lt_axi_s_arcache),
        .i_aic_6_init_lt_axi_s_arid(i_aic_6_init_lt_axi_s_arid),
        .i_aic_6_init_lt_axi_s_arlen(i_aic_6_init_lt_axi_s_arlen),
        .i_aic_6_init_lt_axi_s_arlock(i_aic_6_init_lt_axi_s_arlock),
        .i_aic_6_init_lt_axi_s_arprot(i_aic_6_init_lt_axi_s_arprot),
        .i_aic_6_init_lt_axi_s_arqos(i_aic_6_init_lt_axi_s_arqos),
        .o_aic_6_init_lt_axi_s_arready(o_aic_6_init_lt_axi_s_arready),
        .i_aic_6_init_lt_axi_s_arsize(i_aic_6_init_lt_axi_s_arsize),
        .i_aic_6_init_lt_axi_s_arvalid(i_aic_6_init_lt_axi_s_arvalid),
        .i_aic_6_init_lt_axi_s_awaddr(i_aic_6_init_lt_axi_s_awaddr),
        .i_aic_6_init_lt_axi_s_awburst(i_aic_6_init_lt_axi_s_awburst),
        .i_aic_6_init_lt_axi_s_awcache(i_aic_6_init_lt_axi_s_awcache),
        .i_aic_6_init_lt_axi_s_awid(i_aic_6_init_lt_axi_s_awid),
        .i_aic_6_init_lt_axi_s_awlen(i_aic_6_init_lt_axi_s_awlen),
        .i_aic_6_init_lt_axi_s_awlock(i_aic_6_init_lt_axi_s_awlock),
        .i_aic_6_init_lt_axi_s_awprot(i_aic_6_init_lt_axi_s_awprot),
        .i_aic_6_init_lt_axi_s_awqos(i_aic_6_init_lt_axi_s_awqos),
        .o_aic_6_init_lt_axi_s_awready(o_aic_6_init_lt_axi_s_awready),
        .i_aic_6_init_lt_axi_s_awsize(i_aic_6_init_lt_axi_s_awsize),
        .i_aic_6_init_lt_axi_s_awvalid(i_aic_6_init_lt_axi_s_awvalid),
        .o_aic_6_init_lt_axi_s_bid(o_aic_6_init_lt_axi_s_bid),
        .i_aic_6_init_lt_axi_s_bready(i_aic_6_init_lt_axi_s_bready),
        .o_aic_6_init_lt_axi_s_bresp(o_aic_6_init_lt_axi_s_bresp),
        .o_aic_6_init_lt_axi_s_bvalid(o_aic_6_init_lt_axi_s_bvalid),
        .o_aic_6_init_lt_axi_s_rdata(o_aic_6_init_lt_axi_s_rdata),
        .o_aic_6_init_lt_axi_s_rid(o_aic_6_init_lt_axi_s_rid),
        .o_aic_6_init_lt_axi_s_rlast(o_aic_6_init_lt_axi_s_rlast),
        .i_aic_6_init_lt_axi_s_rready(i_aic_6_init_lt_axi_s_rready),
        .o_aic_6_init_lt_axi_s_rresp(o_aic_6_init_lt_axi_s_rresp),
        .o_aic_6_init_lt_axi_s_rvalid(o_aic_6_init_lt_axi_s_rvalid),
        .i_aic_6_init_lt_axi_s_wdata(i_aic_6_init_lt_axi_s_wdata),
        .i_aic_6_init_lt_axi_s_wlast(i_aic_6_init_lt_axi_s_wlast),
        .o_aic_6_init_lt_axi_s_wready(o_aic_6_init_lt_axi_s_wready),
        .i_aic_6_init_lt_axi_s_wstrb(i_aic_6_init_lt_axi_s_wstrb),
        .i_aic_6_init_lt_axi_s_wvalid(i_aic_6_init_lt_axi_s_wvalid),
        .o_aic_6_pwr_idle_val(o_aic_6_pwr_idle_val),
        .o_aic_6_pwr_idle_ack(o_aic_6_pwr_idle_ack),
        .i_aic_6_pwr_idle_req(i_aic_6_pwr_idle_req),
        .i_aic_6_rst_n(i_aic_6_rst_n),
        .o_aic_6_targ_lt_axi_m_araddr(o_aic_6_targ_lt_axi_m_araddr),
        .o_aic_6_targ_lt_axi_m_arburst(o_aic_6_targ_lt_axi_m_arburst),
        .o_aic_6_targ_lt_axi_m_arcache(o_aic_6_targ_lt_axi_m_arcache),
        .o_aic_6_targ_lt_axi_m_arid(o_aic_6_targ_lt_axi_m_arid),
        .o_aic_6_targ_lt_axi_m_arlen(o_aic_6_targ_lt_axi_m_arlen),
        .o_aic_6_targ_lt_axi_m_arlock(o_aic_6_targ_lt_axi_m_arlock),
        .o_aic_6_targ_lt_axi_m_arprot(o_aic_6_targ_lt_axi_m_arprot),
        .o_aic_6_targ_lt_axi_m_arqos(o_aic_6_targ_lt_axi_m_arqos),
        .i_aic_6_targ_lt_axi_m_arready(i_aic_6_targ_lt_axi_m_arready),
        .o_aic_6_targ_lt_axi_m_arsize(o_aic_6_targ_lt_axi_m_arsize),
        .o_aic_6_targ_lt_axi_m_arvalid(o_aic_6_targ_lt_axi_m_arvalid),
        .o_aic_6_targ_lt_axi_m_awaddr(o_aic_6_targ_lt_axi_m_awaddr),
        .o_aic_6_targ_lt_axi_m_awburst(o_aic_6_targ_lt_axi_m_awburst),
        .o_aic_6_targ_lt_axi_m_awcache(o_aic_6_targ_lt_axi_m_awcache),
        .o_aic_6_targ_lt_axi_m_awid(o_aic_6_targ_lt_axi_m_awid),
        .o_aic_6_targ_lt_axi_m_awlen(o_aic_6_targ_lt_axi_m_awlen),
        .o_aic_6_targ_lt_axi_m_awlock(o_aic_6_targ_lt_axi_m_awlock),
        .o_aic_6_targ_lt_axi_m_awprot(o_aic_6_targ_lt_axi_m_awprot),
        .o_aic_6_targ_lt_axi_m_awqos(o_aic_6_targ_lt_axi_m_awqos),
        .i_aic_6_targ_lt_axi_m_awready(i_aic_6_targ_lt_axi_m_awready),
        .o_aic_6_targ_lt_axi_m_awsize(o_aic_6_targ_lt_axi_m_awsize),
        .o_aic_6_targ_lt_axi_m_awvalid(o_aic_6_targ_lt_axi_m_awvalid),
        .i_aic_6_targ_lt_axi_m_bid(i_aic_6_targ_lt_axi_m_bid),
        .o_aic_6_targ_lt_axi_m_bready(o_aic_6_targ_lt_axi_m_bready),
        .i_aic_6_targ_lt_axi_m_bresp(i_aic_6_targ_lt_axi_m_bresp),
        .i_aic_6_targ_lt_axi_m_bvalid(i_aic_6_targ_lt_axi_m_bvalid),
        .i_aic_6_targ_lt_axi_m_rdata(i_aic_6_targ_lt_axi_m_rdata),
        .i_aic_6_targ_lt_axi_m_rid(i_aic_6_targ_lt_axi_m_rid),
        .i_aic_6_targ_lt_axi_m_rlast(i_aic_6_targ_lt_axi_m_rlast),
        .o_aic_6_targ_lt_axi_m_rready(o_aic_6_targ_lt_axi_m_rready),
        .i_aic_6_targ_lt_axi_m_rresp(i_aic_6_targ_lt_axi_m_rresp),
        .i_aic_6_targ_lt_axi_m_rvalid(i_aic_6_targ_lt_axi_m_rvalid),
        .o_aic_6_targ_lt_axi_m_wdata(o_aic_6_targ_lt_axi_m_wdata),
        .o_aic_6_targ_lt_axi_m_wlast(o_aic_6_targ_lt_axi_m_wlast),
        .i_aic_6_targ_lt_axi_m_wready(i_aic_6_targ_lt_axi_m_wready),
        .o_aic_6_targ_lt_axi_m_wstrb(o_aic_6_targ_lt_axi_m_wstrb),
        .o_aic_6_targ_lt_axi_m_wvalid(o_aic_6_targ_lt_axi_m_wvalid),
        .o_aic_6_targ_syscfg_apb_m_paddr(o_aic_6_targ_syscfg_apb_m_paddr),
        .o_aic_6_targ_syscfg_apb_m_penable(o_aic_6_targ_syscfg_apb_m_penable),
        .o_aic_6_targ_syscfg_apb_m_pprot(o_aic_6_targ_syscfg_apb_m_pprot),
        .i_aic_6_targ_syscfg_apb_m_prdata(i_aic_6_targ_syscfg_apb_m_prdata),
        .i_aic_6_targ_syscfg_apb_m_pready(i_aic_6_targ_syscfg_apb_m_pready),
        .o_aic_6_targ_syscfg_apb_m_psel(o_aic_6_targ_syscfg_apb_m_psel),
        .i_aic_6_targ_syscfg_apb_m_pslverr(i_aic_6_targ_syscfg_apb_m_pslverr),
        .o_aic_6_targ_syscfg_apb_m_pstrb(o_aic_6_targ_syscfg_apb_m_pstrb),
        .o_aic_6_targ_syscfg_apb_m_pwdata(o_aic_6_targ_syscfg_apb_m_pwdata),
        .o_aic_6_targ_syscfg_apb_m_pwrite(o_aic_6_targ_syscfg_apb_m_pwrite),
        .i_aic_7_aon_clk(i_aic_7_aon_clk),
        .i_aic_7_aon_rst_n(i_aic_7_aon_rst_n),
        .i_aic_7_clk(i_aic_7_clk),
        .i_aic_7_clken(i_aic_7_clken),
        .i_aic_7_init_ht_axi_s_araddr(i_aic_7_init_ht_axi_s_araddr),
        .i_aic_7_init_ht_axi_s_arburst(i_aic_7_init_ht_axi_s_arburst),
        .i_aic_7_init_ht_axi_s_arcache(i_aic_7_init_ht_axi_s_arcache),
        .i_aic_7_init_ht_axi_s_arid(i_aic_7_init_ht_axi_s_arid),
        .i_aic_7_init_ht_axi_s_arlen(i_aic_7_init_ht_axi_s_arlen),
        .i_aic_7_init_ht_axi_s_arlock(i_aic_7_init_ht_axi_s_arlock),
        .i_aic_7_init_ht_axi_s_arprot(i_aic_7_init_ht_axi_s_arprot),
        .o_aic_7_init_ht_axi_s_arready(o_aic_7_init_ht_axi_s_arready),
        .i_aic_7_init_ht_axi_s_arsize(i_aic_7_init_ht_axi_s_arsize),
        .i_aic_7_init_ht_axi_s_arvalid(i_aic_7_init_ht_axi_s_arvalid),
        .o_aic_7_init_ht_axi_s_rdata(o_aic_7_init_ht_axi_s_rdata),
        .o_aic_7_init_ht_axi_s_rid(o_aic_7_init_ht_axi_s_rid),
        .o_aic_7_init_ht_axi_s_rlast(o_aic_7_init_ht_axi_s_rlast),
        .i_aic_7_init_ht_axi_s_rready(i_aic_7_init_ht_axi_s_rready),
        .o_aic_7_init_ht_axi_s_rresp(o_aic_7_init_ht_axi_s_rresp),
        .o_aic_7_init_ht_axi_s_rvalid(o_aic_7_init_ht_axi_s_rvalid),
        .i_aic_7_init_ht_axi_s_awaddr(i_aic_7_init_ht_axi_s_awaddr),
        .i_aic_7_init_ht_axi_s_awburst(i_aic_7_init_ht_axi_s_awburst),
        .i_aic_7_init_ht_axi_s_awcache(i_aic_7_init_ht_axi_s_awcache),
        .i_aic_7_init_ht_axi_s_awid(i_aic_7_init_ht_axi_s_awid),
        .i_aic_7_init_ht_axi_s_awlen(i_aic_7_init_ht_axi_s_awlen),
        .i_aic_7_init_ht_axi_s_awlock(i_aic_7_init_ht_axi_s_awlock),
        .i_aic_7_init_ht_axi_s_awprot(i_aic_7_init_ht_axi_s_awprot),
        .o_aic_7_init_ht_axi_s_awready(o_aic_7_init_ht_axi_s_awready),
        .i_aic_7_init_ht_axi_s_awsize(i_aic_7_init_ht_axi_s_awsize),
        .i_aic_7_init_ht_axi_s_awvalid(i_aic_7_init_ht_axi_s_awvalid),
        .o_aic_7_init_ht_axi_s_bid(o_aic_7_init_ht_axi_s_bid),
        .i_aic_7_init_ht_axi_s_bready(i_aic_7_init_ht_axi_s_bready),
        .o_aic_7_init_ht_axi_s_bresp(o_aic_7_init_ht_axi_s_bresp),
        .o_aic_7_init_ht_axi_s_bvalid(o_aic_7_init_ht_axi_s_bvalid),
        .i_aic_7_init_ht_axi_s_wdata(i_aic_7_init_ht_axi_s_wdata),
        .i_aic_7_init_ht_axi_s_wlast(i_aic_7_init_ht_axi_s_wlast),
        .o_aic_7_init_ht_axi_s_wready(o_aic_7_init_ht_axi_s_wready),
        .i_aic_7_init_ht_axi_s_wstrb(i_aic_7_init_ht_axi_s_wstrb),
        .i_aic_7_init_ht_axi_s_wvalid(i_aic_7_init_ht_axi_s_wvalid),
        .i_aic_7_init_lt_axi_s_araddr(i_aic_7_init_lt_axi_s_araddr),
        .i_aic_7_init_lt_axi_s_arburst(i_aic_7_init_lt_axi_s_arburst),
        .i_aic_7_init_lt_axi_s_arcache(i_aic_7_init_lt_axi_s_arcache),
        .i_aic_7_init_lt_axi_s_arid(i_aic_7_init_lt_axi_s_arid),
        .i_aic_7_init_lt_axi_s_arlen(i_aic_7_init_lt_axi_s_arlen),
        .i_aic_7_init_lt_axi_s_arlock(i_aic_7_init_lt_axi_s_arlock),
        .i_aic_7_init_lt_axi_s_arprot(i_aic_7_init_lt_axi_s_arprot),
        .i_aic_7_init_lt_axi_s_arqos(i_aic_7_init_lt_axi_s_arqos),
        .o_aic_7_init_lt_axi_s_arready(o_aic_7_init_lt_axi_s_arready),
        .i_aic_7_init_lt_axi_s_arsize(i_aic_7_init_lt_axi_s_arsize),
        .i_aic_7_init_lt_axi_s_arvalid(i_aic_7_init_lt_axi_s_arvalid),
        .i_aic_7_init_lt_axi_s_awaddr(i_aic_7_init_lt_axi_s_awaddr),
        .i_aic_7_init_lt_axi_s_awburst(i_aic_7_init_lt_axi_s_awburst),
        .i_aic_7_init_lt_axi_s_awcache(i_aic_7_init_lt_axi_s_awcache),
        .i_aic_7_init_lt_axi_s_awid(i_aic_7_init_lt_axi_s_awid),
        .i_aic_7_init_lt_axi_s_awlen(i_aic_7_init_lt_axi_s_awlen),
        .i_aic_7_init_lt_axi_s_awlock(i_aic_7_init_lt_axi_s_awlock),
        .i_aic_7_init_lt_axi_s_awprot(i_aic_7_init_lt_axi_s_awprot),
        .i_aic_7_init_lt_axi_s_awqos(i_aic_7_init_lt_axi_s_awqos),
        .o_aic_7_init_lt_axi_s_awready(o_aic_7_init_lt_axi_s_awready),
        .i_aic_7_init_lt_axi_s_awsize(i_aic_7_init_lt_axi_s_awsize),
        .i_aic_7_init_lt_axi_s_awvalid(i_aic_7_init_lt_axi_s_awvalid),
        .o_aic_7_init_lt_axi_s_bid(o_aic_7_init_lt_axi_s_bid),
        .i_aic_7_init_lt_axi_s_bready(i_aic_7_init_lt_axi_s_bready),
        .o_aic_7_init_lt_axi_s_bresp(o_aic_7_init_lt_axi_s_bresp),
        .o_aic_7_init_lt_axi_s_bvalid(o_aic_7_init_lt_axi_s_bvalid),
        .o_aic_7_init_lt_axi_s_rdata(o_aic_7_init_lt_axi_s_rdata),
        .o_aic_7_init_lt_axi_s_rid(o_aic_7_init_lt_axi_s_rid),
        .o_aic_7_init_lt_axi_s_rlast(o_aic_7_init_lt_axi_s_rlast),
        .i_aic_7_init_lt_axi_s_rready(i_aic_7_init_lt_axi_s_rready),
        .o_aic_7_init_lt_axi_s_rresp(o_aic_7_init_lt_axi_s_rresp),
        .o_aic_7_init_lt_axi_s_rvalid(o_aic_7_init_lt_axi_s_rvalid),
        .i_aic_7_init_lt_axi_s_wdata(i_aic_7_init_lt_axi_s_wdata),
        .i_aic_7_init_lt_axi_s_wlast(i_aic_7_init_lt_axi_s_wlast),
        .o_aic_7_init_lt_axi_s_wready(o_aic_7_init_lt_axi_s_wready),
        .i_aic_7_init_lt_axi_s_wstrb(i_aic_7_init_lt_axi_s_wstrb),
        .i_aic_7_init_lt_axi_s_wvalid(i_aic_7_init_lt_axi_s_wvalid),
        .o_aic_7_pwr_idle_val(o_aic_7_pwr_idle_val),
        .o_aic_7_pwr_idle_ack(o_aic_7_pwr_idle_ack),
        .i_aic_7_pwr_idle_req(i_aic_7_pwr_idle_req),
        .i_aic_7_rst_n(i_aic_7_rst_n),
        .o_aic_7_targ_lt_axi_m_araddr(o_aic_7_targ_lt_axi_m_araddr),
        .o_aic_7_targ_lt_axi_m_arburst(o_aic_7_targ_lt_axi_m_arburst),
        .o_aic_7_targ_lt_axi_m_arcache(o_aic_7_targ_lt_axi_m_arcache),
        .o_aic_7_targ_lt_axi_m_arid(o_aic_7_targ_lt_axi_m_arid),
        .o_aic_7_targ_lt_axi_m_arlen(o_aic_7_targ_lt_axi_m_arlen),
        .o_aic_7_targ_lt_axi_m_arlock(o_aic_7_targ_lt_axi_m_arlock),
        .o_aic_7_targ_lt_axi_m_arprot(o_aic_7_targ_lt_axi_m_arprot),
        .o_aic_7_targ_lt_axi_m_arqos(o_aic_7_targ_lt_axi_m_arqos),
        .i_aic_7_targ_lt_axi_m_arready(i_aic_7_targ_lt_axi_m_arready),
        .o_aic_7_targ_lt_axi_m_arsize(o_aic_7_targ_lt_axi_m_arsize),
        .o_aic_7_targ_lt_axi_m_arvalid(o_aic_7_targ_lt_axi_m_arvalid),
        .o_aic_7_targ_lt_axi_m_awaddr(o_aic_7_targ_lt_axi_m_awaddr),
        .o_aic_7_targ_lt_axi_m_awburst(o_aic_7_targ_lt_axi_m_awburst),
        .o_aic_7_targ_lt_axi_m_awcache(o_aic_7_targ_lt_axi_m_awcache),
        .o_aic_7_targ_lt_axi_m_awid(o_aic_7_targ_lt_axi_m_awid),
        .o_aic_7_targ_lt_axi_m_awlen(o_aic_7_targ_lt_axi_m_awlen),
        .o_aic_7_targ_lt_axi_m_awlock(o_aic_7_targ_lt_axi_m_awlock),
        .o_aic_7_targ_lt_axi_m_awprot(o_aic_7_targ_lt_axi_m_awprot),
        .o_aic_7_targ_lt_axi_m_awqos(o_aic_7_targ_lt_axi_m_awqos),
        .i_aic_7_targ_lt_axi_m_awready(i_aic_7_targ_lt_axi_m_awready),
        .o_aic_7_targ_lt_axi_m_awsize(o_aic_7_targ_lt_axi_m_awsize),
        .o_aic_7_targ_lt_axi_m_awvalid(o_aic_7_targ_lt_axi_m_awvalid),
        .i_aic_7_targ_lt_axi_m_bid(i_aic_7_targ_lt_axi_m_bid),
        .o_aic_7_targ_lt_axi_m_bready(o_aic_7_targ_lt_axi_m_bready),
        .i_aic_7_targ_lt_axi_m_bresp(i_aic_7_targ_lt_axi_m_bresp),
        .i_aic_7_targ_lt_axi_m_bvalid(i_aic_7_targ_lt_axi_m_bvalid),
        .i_aic_7_targ_lt_axi_m_rdata(i_aic_7_targ_lt_axi_m_rdata),
        .i_aic_7_targ_lt_axi_m_rid(i_aic_7_targ_lt_axi_m_rid),
        .i_aic_7_targ_lt_axi_m_rlast(i_aic_7_targ_lt_axi_m_rlast),
        .o_aic_7_targ_lt_axi_m_rready(o_aic_7_targ_lt_axi_m_rready),
        .i_aic_7_targ_lt_axi_m_rresp(i_aic_7_targ_lt_axi_m_rresp),
        .i_aic_7_targ_lt_axi_m_rvalid(i_aic_7_targ_lt_axi_m_rvalid),
        .o_aic_7_targ_lt_axi_m_wdata(o_aic_7_targ_lt_axi_m_wdata),
        .o_aic_7_targ_lt_axi_m_wlast(o_aic_7_targ_lt_axi_m_wlast),
        .i_aic_7_targ_lt_axi_m_wready(i_aic_7_targ_lt_axi_m_wready),
        .o_aic_7_targ_lt_axi_m_wstrb(o_aic_7_targ_lt_axi_m_wstrb),
        .o_aic_7_targ_lt_axi_m_wvalid(o_aic_7_targ_lt_axi_m_wvalid),
        .o_aic_7_targ_syscfg_apb_m_paddr(o_aic_7_targ_syscfg_apb_m_paddr),
        .o_aic_7_targ_syscfg_apb_m_penable(o_aic_7_targ_syscfg_apb_m_penable),
        .o_aic_7_targ_syscfg_apb_m_pprot(o_aic_7_targ_syscfg_apb_m_pprot),
        .i_aic_7_targ_syscfg_apb_m_prdata(i_aic_7_targ_syscfg_apb_m_prdata),
        .i_aic_7_targ_syscfg_apb_m_pready(i_aic_7_targ_syscfg_apb_m_pready),
        .o_aic_7_targ_syscfg_apb_m_psel(o_aic_7_targ_syscfg_apb_m_psel),
        .i_aic_7_targ_syscfg_apb_m_pslverr(i_aic_7_targ_syscfg_apb_m_pslverr),
        .o_aic_7_targ_syscfg_apb_m_pstrb(o_aic_7_targ_syscfg_apb_m_pstrb),
        .o_aic_7_targ_syscfg_apb_m_pwdata(o_aic_7_targ_syscfg_apb_m_pwdata),
        .o_aic_7_targ_syscfg_apb_m_pwrite(o_aic_7_targ_syscfg_apb_m_pwrite),
        .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data),
        .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head),
        .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy),
        .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail),
        .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld),
        .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data),
        .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head),
        .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail),
        .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data),
        .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head),
        .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail),
        .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld),
        .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data),
        .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head),
        .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail),
        .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld),
        .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data),
        .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head),
        .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail),
        .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld),
        .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data),
        .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head),
        .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail),
        .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld),
        .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data),
        .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head),
        .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail),
        .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld),
        .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data),
        .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head),
        .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail),
        .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld),
        .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data),
        .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head),
        .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail),
        .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld),
        .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data),
        .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head),
        .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail),
        .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld),
        .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data),
        .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head),
        .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail),
        .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld),
        .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data),
        .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head),
        .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail),
        .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld),
        .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data),
        .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head),
        .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail),
        .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld),
        .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data),
        .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head),
        .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy),
        .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail),
        .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld),
        .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data),
        .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head),
        .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data),
        .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head),
        .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy),
        .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail),
        .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld),
        .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data),
        .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head),
        .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail),
        .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld),
        .i_l2_4_aon_clk(i_l2_4_aon_clk),
        .i_l2_4_aon_rst_n(i_l2_4_aon_rst_n),
        .i_l2_4_clk(i_l2_4_clk),
        .i_l2_4_clken(i_l2_4_clken),
        .o_l2_4_pwr_idle_val(o_l2_4_pwr_idle_val),
        .o_l2_4_pwr_idle_ack(o_l2_4_pwr_idle_ack),
        .i_l2_4_pwr_idle_req(i_l2_4_pwr_idle_req),
        .i_l2_4_rst_n(i_l2_4_rst_n),
        .o_l2_4_targ_ht_axi_m_araddr(o_l2_4_targ_ht_axi_m_araddr),
        .o_l2_4_targ_ht_axi_m_arburst(o_l2_4_targ_ht_axi_m_arburst),
        .o_l2_4_targ_ht_axi_m_arcache(o_l2_4_targ_ht_axi_m_arcache),
        .o_l2_4_targ_ht_axi_m_arid(o_l2_4_targ_ht_axi_m_arid),
        .o_l2_4_targ_ht_axi_m_arlen(o_l2_4_targ_ht_axi_m_arlen),
        .o_l2_4_targ_ht_axi_m_arlock(o_l2_4_targ_ht_axi_m_arlock),
        .o_l2_4_targ_ht_axi_m_arprot(o_l2_4_targ_ht_axi_m_arprot),
        .i_l2_4_targ_ht_axi_m_arready(i_l2_4_targ_ht_axi_m_arready),
        .o_l2_4_targ_ht_axi_m_arsize(o_l2_4_targ_ht_axi_m_arsize),
        .o_l2_4_targ_ht_axi_m_arvalid(o_l2_4_targ_ht_axi_m_arvalid),
        .i_l2_4_targ_ht_axi_m_rdata(i_l2_4_targ_ht_axi_m_rdata),
        .i_l2_4_targ_ht_axi_m_rid(i_l2_4_targ_ht_axi_m_rid),
        .i_l2_4_targ_ht_axi_m_rlast(i_l2_4_targ_ht_axi_m_rlast),
        .o_l2_4_targ_ht_axi_m_rready(o_l2_4_targ_ht_axi_m_rready),
        .i_l2_4_targ_ht_axi_m_rresp(i_l2_4_targ_ht_axi_m_rresp),
        .i_l2_4_targ_ht_axi_m_rvalid(i_l2_4_targ_ht_axi_m_rvalid),
        .o_l2_4_targ_ht_axi_m_awaddr(o_l2_4_targ_ht_axi_m_awaddr),
        .o_l2_4_targ_ht_axi_m_awburst(o_l2_4_targ_ht_axi_m_awburst),
        .o_l2_4_targ_ht_axi_m_awcache(o_l2_4_targ_ht_axi_m_awcache),
        .o_l2_4_targ_ht_axi_m_awid(o_l2_4_targ_ht_axi_m_awid),
        .o_l2_4_targ_ht_axi_m_awlen(o_l2_4_targ_ht_axi_m_awlen),
        .o_l2_4_targ_ht_axi_m_awlock(o_l2_4_targ_ht_axi_m_awlock),
        .o_l2_4_targ_ht_axi_m_awprot(o_l2_4_targ_ht_axi_m_awprot),
        .i_l2_4_targ_ht_axi_m_awready(i_l2_4_targ_ht_axi_m_awready),
        .o_l2_4_targ_ht_axi_m_awsize(o_l2_4_targ_ht_axi_m_awsize),
        .o_l2_4_targ_ht_axi_m_awvalid(o_l2_4_targ_ht_axi_m_awvalid),
        .i_l2_4_targ_ht_axi_m_bid(i_l2_4_targ_ht_axi_m_bid),
        .o_l2_4_targ_ht_axi_m_bready(o_l2_4_targ_ht_axi_m_bready),
        .i_l2_4_targ_ht_axi_m_bresp(i_l2_4_targ_ht_axi_m_bresp),
        .i_l2_4_targ_ht_axi_m_bvalid(i_l2_4_targ_ht_axi_m_bvalid),
        .o_l2_4_targ_ht_axi_m_wdata(o_l2_4_targ_ht_axi_m_wdata),
        .o_l2_4_targ_ht_axi_m_wlast(o_l2_4_targ_ht_axi_m_wlast),
        .i_l2_4_targ_ht_axi_m_wready(i_l2_4_targ_ht_axi_m_wready),
        .o_l2_4_targ_ht_axi_m_wstrb(o_l2_4_targ_ht_axi_m_wstrb),
        .o_l2_4_targ_ht_axi_m_wvalid(o_l2_4_targ_ht_axi_m_wvalid),
        .o_l2_4_targ_syscfg_apb_m_paddr(o_l2_4_targ_syscfg_apb_m_paddr),
        .o_l2_4_targ_syscfg_apb_m_penable(o_l2_4_targ_syscfg_apb_m_penable),
        .o_l2_4_targ_syscfg_apb_m_pprot(o_l2_4_targ_syscfg_apb_m_pprot),
        .i_l2_4_targ_syscfg_apb_m_prdata(i_l2_4_targ_syscfg_apb_m_prdata),
        .i_l2_4_targ_syscfg_apb_m_pready(i_l2_4_targ_syscfg_apb_m_pready),
        .o_l2_4_targ_syscfg_apb_m_psel(o_l2_4_targ_syscfg_apb_m_psel),
        .i_l2_4_targ_syscfg_apb_m_pslverr(i_l2_4_targ_syscfg_apb_m_pslverr),
        .o_l2_4_targ_syscfg_apb_m_pstrb(o_l2_4_targ_syscfg_apb_m_pstrb),
        .o_l2_4_targ_syscfg_apb_m_pwdata(o_l2_4_targ_syscfg_apb_m_pwdata),
        .o_l2_4_targ_syscfg_apb_m_pwrite(o_l2_4_targ_syscfg_apb_m_pwrite),
        .i_l2_5_aon_clk(i_l2_5_aon_clk),
        .i_l2_5_aon_rst_n(i_l2_5_aon_rst_n),
        .i_l2_5_clk(i_l2_5_clk),
        .i_l2_5_clken(i_l2_5_clken),
        .o_l2_5_pwr_idle_val(o_l2_5_pwr_idle_val),
        .o_l2_5_pwr_idle_ack(o_l2_5_pwr_idle_ack),
        .i_l2_5_pwr_idle_req(i_l2_5_pwr_idle_req),
        .i_l2_5_rst_n(i_l2_5_rst_n),
        .o_l2_5_targ_ht_axi_m_araddr(o_l2_5_targ_ht_axi_m_araddr),
        .o_l2_5_targ_ht_axi_m_arburst(o_l2_5_targ_ht_axi_m_arburst),
        .o_l2_5_targ_ht_axi_m_arcache(o_l2_5_targ_ht_axi_m_arcache),
        .o_l2_5_targ_ht_axi_m_arid(o_l2_5_targ_ht_axi_m_arid),
        .o_l2_5_targ_ht_axi_m_arlen(o_l2_5_targ_ht_axi_m_arlen),
        .o_l2_5_targ_ht_axi_m_arlock(o_l2_5_targ_ht_axi_m_arlock),
        .o_l2_5_targ_ht_axi_m_arprot(o_l2_5_targ_ht_axi_m_arprot),
        .i_l2_5_targ_ht_axi_m_arready(i_l2_5_targ_ht_axi_m_arready),
        .o_l2_5_targ_ht_axi_m_arsize(o_l2_5_targ_ht_axi_m_arsize),
        .o_l2_5_targ_ht_axi_m_arvalid(o_l2_5_targ_ht_axi_m_arvalid),
        .i_l2_5_targ_ht_axi_m_rdata(i_l2_5_targ_ht_axi_m_rdata),
        .i_l2_5_targ_ht_axi_m_rid(i_l2_5_targ_ht_axi_m_rid),
        .i_l2_5_targ_ht_axi_m_rlast(i_l2_5_targ_ht_axi_m_rlast),
        .o_l2_5_targ_ht_axi_m_rready(o_l2_5_targ_ht_axi_m_rready),
        .i_l2_5_targ_ht_axi_m_rresp(i_l2_5_targ_ht_axi_m_rresp),
        .i_l2_5_targ_ht_axi_m_rvalid(i_l2_5_targ_ht_axi_m_rvalid),
        .o_l2_5_targ_ht_axi_m_awaddr(o_l2_5_targ_ht_axi_m_awaddr),
        .o_l2_5_targ_ht_axi_m_awburst(o_l2_5_targ_ht_axi_m_awburst),
        .o_l2_5_targ_ht_axi_m_awcache(o_l2_5_targ_ht_axi_m_awcache),
        .o_l2_5_targ_ht_axi_m_awid(o_l2_5_targ_ht_axi_m_awid),
        .o_l2_5_targ_ht_axi_m_awlen(o_l2_5_targ_ht_axi_m_awlen),
        .o_l2_5_targ_ht_axi_m_awlock(o_l2_5_targ_ht_axi_m_awlock),
        .o_l2_5_targ_ht_axi_m_awprot(o_l2_5_targ_ht_axi_m_awprot),
        .i_l2_5_targ_ht_axi_m_awready(i_l2_5_targ_ht_axi_m_awready),
        .o_l2_5_targ_ht_axi_m_awsize(o_l2_5_targ_ht_axi_m_awsize),
        .o_l2_5_targ_ht_axi_m_awvalid(o_l2_5_targ_ht_axi_m_awvalid),
        .i_l2_5_targ_ht_axi_m_bid(i_l2_5_targ_ht_axi_m_bid),
        .o_l2_5_targ_ht_axi_m_bready(o_l2_5_targ_ht_axi_m_bready),
        .i_l2_5_targ_ht_axi_m_bresp(i_l2_5_targ_ht_axi_m_bresp),
        .i_l2_5_targ_ht_axi_m_bvalid(i_l2_5_targ_ht_axi_m_bvalid),
        .o_l2_5_targ_ht_axi_m_wdata(o_l2_5_targ_ht_axi_m_wdata),
        .o_l2_5_targ_ht_axi_m_wlast(o_l2_5_targ_ht_axi_m_wlast),
        .i_l2_5_targ_ht_axi_m_wready(i_l2_5_targ_ht_axi_m_wready),
        .o_l2_5_targ_ht_axi_m_wstrb(o_l2_5_targ_ht_axi_m_wstrb),
        .o_l2_5_targ_ht_axi_m_wvalid(o_l2_5_targ_ht_axi_m_wvalid),
        .o_l2_5_targ_syscfg_apb_m_paddr(o_l2_5_targ_syscfg_apb_m_paddr),
        .o_l2_5_targ_syscfg_apb_m_penable(o_l2_5_targ_syscfg_apb_m_penable),
        .o_l2_5_targ_syscfg_apb_m_pprot(o_l2_5_targ_syscfg_apb_m_pprot),
        .i_l2_5_targ_syscfg_apb_m_prdata(i_l2_5_targ_syscfg_apb_m_prdata),
        .i_l2_5_targ_syscfg_apb_m_pready(i_l2_5_targ_syscfg_apb_m_pready),
        .o_l2_5_targ_syscfg_apb_m_psel(o_l2_5_targ_syscfg_apb_m_psel),
        .i_l2_5_targ_syscfg_apb_m_pslverr(i_l2_5_targ_syscfg_apb_m_pslverr),
        .o_l2_5_targ_syscfg_apb_m_pstrb(o_l2_5_targ_syscfg_apb_m_pstrb),
        .o_l2_5_targ_syscfg_apb_m_pwdata(o_l2_5_targ_syscfg_apb_m_pwdata),
        .o_l2_5_targ_syscfg_apb_m_pwrite(o_l2_5_targ_syscfg_apb_m_pwrite),
        .i_l2_6_aon_clk(i_l2_6_aon_clk),
        .i_l2_6_aon_rst_n(i_l2_6_aon_rst_n),
        .i_l2_6_clk(i_l2_6_clk),
        .i_l2_6_clken(i_l2_6_clken),
        .o_l2_6_pwr_idle_val(o_l2_6_pwr_idle_val),
        .o_l2_6_pwr_idle_ack(o_l2_6_pwr_idle_ack),
        .i_l2_6_pwr_idle_req(i_l2_6_pwr_idle_req),
        .i_l2_6_rst_n(i_l2_6_rst_n),
        .o_l2_6_targ_ht_axi_m_araddr(o_l2_6_targ_ht_axi_m_araddr),
        .o_l2_6_targ_ht_axi_m_arburst(o_l2_6_targ_ht_axi_m_arburst),
        .o_l2_6_targ_ht_axi_m_arcache(o_l2_6_targ_ht_axi_m_arcache),
        .o_l2_6_targ_ht_axi_m_arid(o_l2_6_targ_ht_axi_m_arid),
        .o_l2_6_targ_ht_axi_m_arlen(o_l2_6_targ_ht_axi_m_arlen),
        .o_l2_6_targ_ht_axi_m_arlock(o_l2_6_targ_ht_axi_m_arlock),
        .o_l2_6_targ_ht_axi_m_arprot(o_l2_6_targ_ht_axi_m_arprot),
        .i_l2_6_targ_ht_axi_m_arready(i_l2_6_targ_ht_axi_m_arready),
        .o_l2_6_targ_ht_axi_m_arsize(o_l2_6_targ_ht_axi_m_arsize),
        .o_l2_6_targ_ht_axi_m_arvalid(o_l2_6_targ_ht_axi_m_arvalid),
        .i_l2_6_targ_ht_axi_m_rdata(i_l2_6_targ_ht_axi_m_rdata),
        .i_l2_6_targ_ht_axi_m_rid(i_l2_6_targ_ht_axi_m_rid),
        .i_l2_6_targ_ht_axi_m_rlast(i_l2_6_targ_ht_axi_m_rlast),
        .o_l2_6_targ_ht_axi_m_rready(o_l2_6_targ_ht_axi_m_rready),
        .i_l2_6_targ_ht_axi_m_rresp(i_l2_6_targ_ht_axi_m_rresp),
        .i_l2_6_targ_ht_axi_m_rvalid(i_l2_6_targ_ht_axi_m_rvalid),
        .o_l2_6_targ_ht_axi_m_awaddr(o_l2_6_targ_ht_axi_m_awaddr),
        .o_l2_6_targ_ht_axi_m_awburst(o_l2_6_targ_ht_axi_m_awburst),
        .o_l2_6_targ_ht_axi_m_awcache(o_l2_6_targ_ht_axi_m_awcache),
        .o_l2_6_targ_ht_axi_m_awid(o_l2_6_targ_ht_axi_m_awid),
        .o_l2_6_targ_ht_axi_m_awlen(o_l2_6_targ_ht_axi_m_awlen),
        .o_l2_6_targ_ht_axi_m_awlock(o_l2_6_targ_ht_axi_m_awlock),
        .o_l2_6_targ_ht_axi_m_awprot(o_l2_6_targ_ht_axi_m_awprot),
        .i_l2_6_targ_ht_axi_m_awready(i_l2_6_targ_ht_axi_m_awready),
        .o_l2_6_targ_ht_axi_m_awsize(o_l2_6_targ_ht_axi_m_awsize),
        .o_l2_6_targ_ht_axi_m_awvalid(o_l2_6_targ_ht_axi_m_awvalid),
        .i_l2_6_targ_ht_axi_m_bid(i_l2_6_targ_ht_axi_m_bid),
        .o_l2_6_targ_ht_axi_m_bready(o_l2_6_targ_ht_axi_m_bready),
        .i_l2_6_targ_ht_axi_m_bresp(i_l2_6_targ_ht_axi_m_bresp),
        .i_l2_6_targ_ht_axi_m_bvalid(i_l2_6_targ_ht_axi_m_bvalid),
        .o_l2_6_targ_ht_axi_m_wdata(o_l2_6_targ_ht_axi_m_wdata),
        .o_l2_6_targ_ht_axi_m_wlast(o_l2_6_targ_ht_axi_m_wlast),
        .i_l2_6_targ_ht_axi_m_wready(i_l2_6_targ_ht_axi_m_wready),
        .o_l2_6_targ_ht_axi_m_wstrb(o_l2_6_targ_ht_axi_m_wstrb),
        .o_l2_6_targ_ht_axi_m_wvalid(o_l2_6_targ_ht_axi_m_wvalid),
        .o_l2_6_targ_syscfg_apb_m_paddr(o_l2_6_targ_syscfg_apb_m_paddr),
        .o_l2_6_targ_syscfg_apb_m_penable(o_l2_6_targ_syscfg_apb_m_penable),
        .o_l2_6_targ_syscfg_apb_m_pprot(o_l2_6_targ_syscfg_apb_m_pprot),
        .i_l2_6_targ_syscfg_apb_m_prdata(i_l2_6_targ_syscfg_apb_m_prdata),
        .i_l2_6_targ_syscfg_apb_m_pready(i_l2_6_targ_syscfg_apb_m_pready),
        .o_l2_6_targ_syscfg_apb_m_psel(o_l2_6_targ_syscfg_apb_m_psel),
        .i_l2_6_targ_syscfg_apb_m_pslverr(i_l2_6_targ_syscfg_apb_m_pslverr),
        .o_l2_6_targ_syscfg_apb_m_pstrb(o_l2_6_targ_syscfg_apb_m_pstrb),
        .o_l2_6_targ_syscfg_apb_m_pwdata(o_l2_6_targ_syscfg_apb_m_pwdata),
        .o_l2_6_targ_syscfg_apb_m_pwrite(o_l2_6_targ_syscfg_apb_m_pwrite),
        .i_l2_7_aon_clk(i_l2_7_aon_clk),
        .i_l2_7_aon_rst_n(i_l2_7_aon_rst_n),
        .i_l2_7_clk(i_l2_7_clk),
        .i_l2_7_clken(i_l2_7_clken),
        .o_l2_7_pwr_idle_val(o_l2_7_pwr_idle_val),
        .o_l2_7_pwr_idle_ack(o_l2_7_pwr_idle_ack),
        .i_l2_7_pwr_idle_req(i_l2_7_pwr_idle_req),
        .i_l2_7_rst_n(i_l2_7_rst_n),
        .o_l2_7_targ_ht_axi_m_araddr(o_l2_7_targ_ht_axi_m_araddr),
        .o_l2_7_targ_ht_axi_m_arburst(o_l2_7_targ_ht_axi_m_arburst),
        .o_l2_7_targ_ht_axi_m_arcache(o_l2_7_targ_ht_axi_m_arcache),
        .o_l2_7_targ_ht_axi_m_arid(o_l2_7_targ_ht_axi_m_arid),
        .o_l2_7_targ_ht_axi_m_arlen(o_l2_7_targ_ht_axi_m_arlen),
        .o_l2_7_targ_ht_axi_m_arlock(o_l2_7_targ_ht_axi_m_arlock),
        .o_l2_7_targ_ht_axi_m_arprot(o_l2_7_targ_ht_axi_m_arprot),
        .i_l2_7_targ_ht_axi_m_arready(i_l2_7_targ_ht_axi_m_arready),
        .o_l2_7_targ_ht_axi_m_arsize(o_l2_7_targ_ht_axi_m_arsize),
        .o_l2_7_targ_ht_axi_m_arvalid(o_l2_7_targ_ht_axi_m_arvalid),
        .i_l2_7_targ_ht_axi_m_rdata(i_l2_7_targ_ht_axi_m_rdata),
        .i_l2_7_targ_ht_axi_m_rid(i_l2_7_targ_ht_axi_m_rid),
        .i_l2_7_targ_ht_axi_m_rlast(i_l2_7_targ_ht_axi_m_rlast),
        .o_l2_7_targ_ht_axi_m_rready(o_l2_7_targ_ht_axi_m_rready),
        .i_l2_7_targ_ht_axi_m_rresp(i_l2_7_targ_ht_axi_m_rresp),
        .i_l2_7_targ_ht_axi_m_rvalid(i_l2_7_targ_ht_axi_m_rvalid),
        .o_l2_7_targ_ht_axi_m_awaddr(o_l2_7_targ_ht_axi_m_awaddr),
        .o_l2_7_targ_ht_axi_m_awburst(o_l2_7_targ_ht_axi_m_awburst),
        .o_l2_7_targ_ht_axi_m_awcache(o_l2_7_targ_ht_axi_m_awcache),
        .o_l2_7_targ_ht_axi_m_awid(o_l2_7_targ_ht_axi_m_awid),
        .o_l2_7_targ_ht_axi_m_awlen(o_l2_7_targ_ht_axi_m_awlen),
        .o_l2_7_targ_ht_axi_m_awlock(o_l2_7_targ_ht_axi_m_awlock),
        .o_l2_7_targ_ht_axi_m_awprot(o_l2_7_targ_ht_axi_m_awprot),
        .i_l2_7_targ_ht_axi_m_awready(i_l2_7_targ_ht_axi_m_awready),
        .o_l2_7_targ_ht_axi_m_awsize(o_l2_7_targ_ht_axi_m_awsize),
        .o_l2_7_targ_ht_axi_m_awvalid(o_l2_7_targ_ht_axi_m_awvalid),
        .i_l2_7_targ_ht_axi_m_bid(i_l2_7_targ_ht_axi_m_bid),
        .o_l2_7_targ_ht_axi_m_bready(o_l2_7_targ_ht_axi_m_bready),
        .i_l2_7_targ_ht_axi_m_bresp(i_l2_7_targ_ht_axi_m_bresp),
        .i_l2_7_targ_ht_axi_m_bvalid(i_l2_7_targ_ht_axi_m_bvalid),
        .o_l2_7_targ_ht_axi_m_wdata(o_l2_7_targ_ht_axi_m_wdata),
        .o_l2_7_targ_ht_axi_m_wlast(o_l2_7_targ_ht_axi_m_wlast),
        .i_l2_7_targ_ht_axi_m_wready(i_l2_7_targ_ht_axi_m_wready),
        .o_l2_7_targ_ht_axi_m_wstrb(o_l2_7_targ_ht_axi_m_wstrb),
        .o_l2_7_targ_ht_axi_m_wvalid(o_l2_7_targ_ht_axi_m_wvalid),
        .o_l2_7_targ_syscfg_apb_m_paddr(o_l2_7_targ_syscfg_apb_m_paddr),
        .o_l2_7_targ_syscfg_apb_m_penable(o_l2_7_targ_syscfg_apb_m_penable),
        .o_l2_7_targ_syscfg_apb_m_pprot(o_l2_7_targ_syscfg_apb_m_pprot),
        .i_l2_7_targ_syscfg_apb_m_prdata(i_l2_7_targ_syscfg_apb_m_prdata),
        .i_l2_7_targ_syscfg_apb_m_pready(i_l2_7_targ_syscfg_apb_m_pready),
        .o_l2_7_targ_syscfg_apb_m_psel(o_l2_7_targ_syscfg_apb_m_psel),
        .i_l2_7_targ_syscfg_apb_m_pslverr(i_l2_7_targ_syscfg_apb_m_pslverr),
        .o_l2_7_targ_syscfg_apb_m_pstrb(o_l2_7_targ_syscfg_apb_m_pstrb),
        .o_l2_7_targ_syscfg_apb_m_pwdata(o_l2_7_targ_syscfg_apb_m_pwdata),
        .o_l2_7_targ_syscfg_apb_m_pwrite(o_l2_7_targ_syscfg_apb_m_pwrite),
        .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
        .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
        .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
        .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
        .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
        .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
        .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
        .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
        .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
        .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
        .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
        .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),

        // Token Network IOs
        // - Fences
        .o_aic_4_pwr_tok_idle_val(o_aic_4_pwr_tok_idle_val),
        .o_aic_4_pwr_tok_idle_ack(o_aic_4_pwr_tok_idle_ack),
        .i_aic_4_pwr_tok_idle_req(i_aic_4_pwr_tok_idle_req),
        .o_aic_5_pwr_tok_idle_val(o_aic_5_pwr_tok_idle_val),
        .o_aic_5_pwr_tok_idle_ack(o_aic_5_pwr_tok_idle_ack),
        .i_aic_5_pwr_tok_idle_req(i_aic_5_pwr_tok_idle_req),
        .o_aic_6_pwr_tok_idle_val(o_aic_6_pwr_tok_idle_val),
        .o_aic_6_pwr_tok_idle_ack(o_aic_6_pwr_tok_idle_ack),
        .i_aic_6_pwr_tok_idle_req(i_aic_6_pwr_tok_idle_req),
        .o_aic_7_pwr_tok_idle_val(o_aic_7_pwr_tok_idle_val),
        .o_aic_7_pwr_tok_idle_ack(o_aic_7_pwr_tok_idle_ack),
        .i_aic_7_pwr_tok_idle_req(i_aic_7_pwr_tok_idle_req),

        // - NIUs
        .i_aic_4_init_tok_ocpl_s_maddr     (i_aic_4_init_tok_ocpl_s_maddr),
        .i_aic_4_init_tok_ocpl_s_mcmd      (i_aic_4_init_tok_ocpl_s_mcmd),
        .i_aic_4_init_tok_ocpl_s_mdata     (i_aic_4_init_tok_ocpl_s_mdata),
        .o_aic_4_init_tok_ocpl_s_scmdaccept(o_aic_4_init_tok_ocpl_s_scmdaccept),
        .o_aic_4_targ_tok_ocpl_m_maddr     (o_aic_4_targ_tok_ocpl_m_maddr),
        .o_aic_4_targ_tok_ocpl_m_mcmd      (o_aic_4_targ_tok_ocpl_m_mcmd),
        .o_aic_4_targ_tok_ocpl_m_mdata     (o_aic_4_targ_tok_ocpl_m_mdata),
        .i_aic_4_targ_tok_ocpl_m_scmdaccept(i_aic_4_targ_tok_ocpl_m_scmdaccept),
        .i_aic_5_init_tok_ocpl_s_maddr     (i_aic_5_init_tok_ocpl_s_maddr),
        .i_aic_5_init_tok_ocpl_s_mcmd      (i_aic_5_init_tok_ocpl_s_mcmd),
        .i_aic_5_init_tok_ocpl_s_mdata     (i_aic_5_init_tok_ocpl_s_mdata),
        .o_aic_5_init_tok_ocpl_s_scmdaccept(o_aic_5_init_tok_ocpl_s_scmdaccept),
        .o_aic_5_targ_tok_ocpl_m_maddr     (o_aic_5_targ_tok_ocpl_m_maddr),
        .o_aic_5_targ_tok_ocpl_m_mcmd      (o_aic_5_targ_tok_ocpl_m_mcmd),
        .o_aic_5_targ_tok_ocpl_m_mdata     (o_aic_5_targ_tok_ocpl_m_mdata),
        .i_aic_5_targ_tok_ocpl_m_scmdaccept(i_aic_5_targ_tok_ocpl_m_scmdaccept),
        .i_aic_6_init_tok_ocpl_s_maddr     (i_aic_6_init_tok_ocpl_s_maddr),
        .i_aic_6_init_tok_ocpl_s_mcmd      (i_aic_6_init_tok_ocpl_s_mcmd),
        .i_aic_6_init_tok_ocpl_s_mdata     (i_aic_6_init_tok_ocpl_s_mdata),
        .o_aic_6_init_tok_ocpl_s_scmdaccept(o_aic_6_init_tok_ocpl_s_scmdaccept),
        .o_aic_6_targ_tok_ocpl_m_maddr     (o_aic_6_targ_tok_ocpl_m_maddr),
        .o_aic_6_targ_tok_ocpl_m_mcmd      (o_aic_6_targ_tok_ocpl_m_mcmd),
        .o_aic_6_targ_tok_ocpl_m_mdata     (o_aic_6_targ_tok_ocpl_m_mdata),
        .i_aic_6_targ_tok_ocpl_m_scmdaccept(i_aic_6_targ_tok_ocpl_m_scmdaccept),
        .i_aic_7_init_tok_ocpl_s_maddr     (i_aic_7_init_tok_ocpl_s_maddr),
        .i_aic_7_init_tok_ocpl_s_mcmd      (i_aic_7_init_tok_ocpl_s_mcmd),
        .i_aic_7_init_tok_ocpl_s_mdata     (i_aic_7_init_tok_ocpl_s_mdata),
        .o_aic_7_init_tok_ocpl_s_scmdaccept(o_aic_7_init_tok_ocpl_s_scmdaccept),
        .o_aic_7_targ_tok_ocpl_m_maddr     (o_aic_7_targ_tok_ocpl_m_maddr),
        .o_aic_7_targ_tok_ocpl_m_mcmd      (o_aic_7_targ_tok_ocpl_m_mcmd),
        .o_aic_7_targ_tok_ocpl_m_mdata     (o_aic_7_targ_tok_ocpl_m_mdata),
        .i_aic_7_targ_tok_ocpl_m_scmdaccept(i_aic_7_targ_tok_ocpl_m_scmdaccept),

        .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data),
        .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head),
        .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy),
        .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail),
        .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld),
        .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data),
        .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head),
        .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy),
        .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail),
        .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld),
        .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data),
        .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head),
        .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy),
        .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail),
        .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld),
        .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data),
        .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head),
        .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy),
        .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail),
        .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld),

        .i_noc_clk(i_noc_clk),
        .i_noc_rst_n(i_noc_rst_n),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  )
    );

    // Instance of noc_h_south_p
    noc_h_south_p h_south_p (
        .i_aic_0_aon_clk(i_aic_0_aon_clk),
        .i_aic_0_aon_rst_n(i_aic_0_aon_rst_n),
        .i_aic_0_clk(i_aic_0_clk),
        .i_aic_0_clken(i_aic_0_clken),
        .i_aic_0_init_ht_axi_s_araddr(i_aic_0_init_ht_axi_s_araddr),
        .i_aic_0_init_ht_axi_s_arburst(i_aic_0_init_ht_axi_s_arburst),
        .i_aic_0_init_ht_axi_s_arcache(i_aic_0_init_ht_axi_s_arcache),
        .i_aic_0_init_ht_axi_s_arid(i_aic_0_init_ht_axi_s_arid),
        .i_aic_0_init_ht_axi_s_arlen(i_aic_0_init_ht_axi_s_arlen),
        .i_aic_0_init_ht_axi_s_arlock(i_aic_0_init_ht_axi_s_arlock),
        .i_aic_0_init_ht_axi_s_arprot(i_aic_0_init_ht_axi_s_arprot),
        .o_aic_0_init_ht_axi_s_arready(o_aic_0_init_ht_axi_s_arready),
        .i_aic_0_init_ht_axi_s_arsize(i_aic_0_init_ht_axi_s_arsize),
        .i_aic_0_init_ht_axi_s_arvalid(i_aic_0_init_ht_axi_s_arvalid),
        .o_aic_0_init_ht_axi_s_rdata(o_aic_0_init_ht_axi_s_rdata),
        .o_aic_0_init_ht_axi_s_rid(o_aic_0_init_ht_axi_s_rid),
        .o_aic_0_init_ht_axi_s_rlast(o_aic_0_init_ht_axi_s_rlast),
        .i_aic_0_init_ht_axi_s_rready(i_aic_0_init_ht_axi_s_rready),
        .o_aic_0_init_ht_axi_s_rresp(o_aic_0_init_ht_axi_s_rresp),
        .o_aic_0_init_ht_axi_s_rvalid(o_aic_0_init_ht_axi_s_rvalid),
        .i_aic_0_init_ht_axi_s_awaddr(i_aic_0_init_ht_axi_s_awaddr),
        .i_aic_0_init_ht_axi_s_awburst(i_aic_0_init_ht_axi_s_awburst),
        .i_aic_0_init_ht_axi_s_awcache(i_aic_0_init_ht_axi_s_awcache),
        .i_aic_0_init_ht_axi_s_awid(i_aic_0_init_ht_axi_s_awid),
        .i_aic_0_init_ht_axi_s_awlen(i_aic_0_init_ht_axi_s_awlen),
        .i_aic_0_init_ht_axi_s_awlock(i_aic_0_init_ht_axi_s_awlock),
        .i_aic_0_init_ht_axi_s_awprot(i_aic_0_init_ht_axi_s_awprot),
        .o_aic_0_init_ht_axi_s_awready(o_aic_0_init_ht_axi_s_awready),
        .i_aic_0_init_ht_axi_s_awsize(i_aic_0_init_ht_axi_s_awsize),
        .i_aic_0_init_ht_axi_s_awvalid(i_aic_0_init_ht_axi_s_awvalid),
        .o_aic_0_init_ht_axi_s_bid(o_aic_0_init_ht_axi_s_bid),
        .i_aic_0_init_ht_axi_s_bready(i_aic_0_init_ht_axi_s_bready),
        .o_aic_0_init_ht_axi_s_bresp(o_aic_0_init_ht_axi_s_bresp),
        .o_aic_0_init_ht_axi_s_bvalid(o_aic_0_init_ht_axi_s_bvalid),
        .i_aic_0_init_ht_axi_s_wdata(i_aic_0_init_ht_axi_s_wdata),
        .i_aic_0_init_ht_axi_s_wlast(i_aic_0_init_ht_axi_s_wlast),
        .o_aic_0_init_ht_axi_s_wready(o_aic_0_init_ht_axi_s_wready),
        .i_aic_0_init_ht_axi_s_wstrb(i_aic_0_init_ht_axi_s_wstrb),
        .i_aic_0_init_ht_axi_s_wvalid(i_aic_0_init_ht_axi_s_wvalid),
        .i_aic_0_init_lt_axi_s_araddr(i_aic_0_init_lt_axi_s_araddr),
        .i_aic_0_init_lt_axi_s_arburst(i_aic_0_init_lt_axi_s_arburst),
        .i_aic_0_init_lt_axi_s_arcache(i_aic_0_init_lt_axi_s_arcache),
        .i_aic_0_init_lt_axi_s_arid(i_aic_0_init_lt_axi_s_arid),
        .i_aic_0_init_lt_axi_s_arlen(i_aic_0_init_lt_axi_s_arlen),
        .i_aic_0_init_lt_axi_s_arlock(i_aic_0_init_lt_axi_s_arlock),
        .i_aic_0_init_lt_axi_s_arprot(i_aic_0_init_lt_axi_s_arprot),
        .i_aic_0_init_lt_axi_s_arqos(i_aic_0_init_lt_axi_s_arqos),
        .o_aic_0_init_lt_axi_s_arready(o_aic_0_init_lt_axi_s_arready),
        .i_aic_0_init_lt_axi_s_arsize(i_aic_0_init_lt_axi_s_arsize),
        .i_aic_0_init_lt_axi_s_arvalid(i_aic_0_init_lt_axi_s_arvalid),
        .i_aic_0_init_lt_axi_s_awaddr(i_aic_0_init_lt_axi_s_awaddr),
        .i_aic_0_init_lt_axi_s_awburst(i_aic_0_init_lt_axi_s_awburst),
        .i_aic_0_init_lt_axi_s_awcache(i_aic_0_init_lt_axi_s_awcache),
        .i_aic_0_init_lt_axi_s_awid(i_aic_0_init_lt_axi_s_awid),
        .i_aic_0_init_lt_axi_s_awlen(i_aic_0_init_lt_axi_s_awlen),
        .i_aic_0_init_lt_axi_s_awlock(i_aic_0_init_lt_axi_s_awlock),
        .i_aic_0_init_lt_axi_s_awprot(i_aic_0_init_lt_axi_s_awprot),
        .i_aic_0_init_lt_axi_s_awqos(i_aic_0_init_lt_axi_s_awqos),
        .o_aic_0_init_lt_axi_s_awready(o_aic_0_init_lt_axi_s_awready),
        .i_aic_0_init_lt_axi_s_awsize(i_aic_0_init_lt_axi_s_awsize),
        .i_aic_0_init_lt_axi_s_awvalid(i_aic_0_init_lt_axi_s_awvalid),
        .o_aic_0_init_lt_axi_s_bid(o_aic_0_init_lt_axi_s_bid),
        .i_aic_0_init_lt_axi_s_bready(i_aic_0_init_lt_axi_s_bready),
        .o_aic_0_init_lt_axi_s_bresp(o_aic_0_init_lt_axi_s_bresp),
        .o_aic_0_init_lt_axi_s_bvalid(o_aic_0_init_lt_axi_s_bvalid),
        .o_aic_0_init_lt_axi_s_rdata(o_aic_0_init_lt_axi_s_rdata),
        .o_aic_0_init_lt_axi_s_rid(o_aic_0_init_lt_axi_s_rid),
        .o_aic_0_init_lt_axi_s_rlast(o_aic_0_init_lt_axi_s_rlast),
        .i_aic_0_init_lt_axi_s_rready(i_aic_0_init_lt_axi_s_rready),
        .o_aic_0_init_lt_axi_s_rresp(o_aic_0_init_lt_axi_s_rresp),
        .o_aic_0_init_lt_axi_s_rvalid(o_aic_0_init_lt_axi_s_rvalid),
        .i_aic_0_init_lt_axi_s_wdata(i_aic_0_init_lt_axi_s_wdata),
        .i_aic_0_init_lt_axi_s_wlast(i_aic_0_init_lt_axi_s_wlast),
        .o_aic_0_init_lt_axi_s_wready(o_aic_0_init_lt_axi_s_wready),
        .i_aic_0_init_lt_axi_s_wstrb(i_aic_0_init_lt_axi_s_wstrb),
        .i_aic_0_init_lt_axi_s_wvalid(i_aic_0_init_lt_axi_s_wvalid),
        .o_aic_0_pwr_idle_val(o_aic_0_pwr_idle_val),
        .o_aic_0_pwr_idle_ack(o_aic_0_pwr_idle_ack),
        .i_aic_0_pwr_idle_req(i_aic_0_pwr_idle_req),
        .i_aic_0_rst_n(i_aic_0_rst_n),
        .o_aic_0_targ_lt_axi_m_araddr(o_aic_0_targ_lt_axi_m_araddr),
        .o_aic_0_targ_lt_axi_m_arburst(o_aic_0_targ_lt_axi_m_arburst),
        .o_aic_0_targ_lt_axi_m_arcache(o_aic_0_targ_lt_axi_m_arcache),
        .o_aic_0_targ_lt_axi_m_arid(o_aic_0_targ_lt_axi_m_arid),
        .o_aic_0_targ_lt_axi_m_arlen(o_aic_0_targ_lt_axi_m_arlen),
        .o_aic_0_targ_lt_axi_m_arlock(o_aic_0_targ_lt_axi_m_arlock),
        .o_aic_0_targ_lt_axi_m_arprot(o_aic_0_targ_lt_axi_m_arprot),
        .o_aic_0_targ_lt_axi_m_arqos(o_aic_0_targ_lt_axi_m_arqos),
        .i_aic_0_targ_lt_axi_m_arready(i_aic_0_targ_lt_axi_m_arready),
        .o_aic_0_targ_lt_axi_m_arsize(o_aic_0_targ_lt_axi_m_arsize),
        .o_aic_0_targ_lt_axi_m_arvalid(o_aic_0_targ_lt_axi_m_arvalid),
        .o_aic_0_targ_lt_axi_m_awaddr(o_aic_0_targ_lt_axi_m_awaddr),
        .o_aic_0_targ_lt_axi_m_awburst(o_aic_0_targ_lt_axi_m_awburst),
        .o_aic_0_targ_lt_axi_m_awcache(o_aic_0_targ_lt_axi_m_awcache),
        .o_aic_0_targ_lt_axi_m_awid(o_aic_0_targ_lt_axi_m_awid),
        .o_aic_0_targ_lt_axi_m_awlen(o_aic_0_targ_lt_axi_m_awlen),
        .o_aic_0_targ_lt_axi_m_awlock(o_aic_0_targ_lt_axi_m_awlock),
        .o_aic_0_targ_lt_axi_m_awprot(o_aic_0_targ_lt_axi_m_awprot),
        .o_aic_0_targ_lt_axi_m_awqos(o_aic_0_targ_lt_axi_m_awqos),
        .i_aic_0_targ_lt_axi_m_awready(i_aic_0_targ_lt_axi_m_awready),
        .o_aic_0_targ_lt_axi_m_awsize(o_aic_0_targ_lt_axi_m_awsize),
        .o_aic_0_targ_lt_axi_m_awvalid(o_aic_0_targ_lt_axi_m_awvalid),
        .i_aic_0_targ_lt_axi_m_bid(i_aic_0_targ_lt_axi_m_bid),
        .o_aic_0_targ_lt_axi_m_bready(o_aic_0_targ_lt_axi_m_bready),
        .i_aic_0_targ_lt_axi_m_bresp(i_aic_0_targ_lt_axi_m_bresp),
        .i_aic_0_targ_lt_axi_m_bvalid(i_aic_0_targ_lt_axi_m_bvalid),
        .i_aic_0_targ_lt_axi_m_rdata(i_aic_0_targ_lt_axi_m_rdata),
        .i_aic_0_targ_lt_axi_m_rid(i_aic_0_targ_lt_axi_m_rid),
        .i_aic_0_targ_lt_axi_m_rlast(i_aic_0_targ_lt_axi_m_rlast),
        .o_aic_0_targ_lt_axi_m_rready(o_aic_0_targ_lt_axi_m_rready),
        .i_aic_0_targ_lt_axi_m_rresp(i_aic_0_targ_lt_axi_m_rresp),
        .i_aic_0_targ_lt_axi_m_rvalid(i_aic_0_targ_lt_axi_m_rvalid),
        .o_aic_0_targ_lt_axi_m_wdata(o_aic_0_targ_lt_axi_m_wdata),
        .o_aic_0_targ_lt_axi_m_wlast(o_aic_0_targ_lt_axi_m_wlast),
        .i_aic_0_targ_lt_axi_m_wready(i_aic_0_targ_lt_axi_m_wready),
        .o_aic_0_targ_lt_axi_m_wstrb(o_aic_0_targ_lt_axi_m_wstrb),
        .o_aic_0_targ_lt_axi_m_wvalid(o_aic_0_targ_lt_axi_m_wvalid),
        .o_aic_0_targ_syscfg_apb_m_paddr(o_aic_0_targ_syscfg_apb_m_paddr),
        .o_aic_0_targ_syscfg_apb_m_penable(o_aic_0_targ_syscfg_apb_m_penable),
        .o_aic_0_targ_syscfg_apb_m_pprot(o_aic_0_targ_syscfg_apb_m_pprot),
        .i_aic_0_targ_syscfg_apb_m_prdata(i_aic_0_targ_syscfg_apb_m_prdata),
        .i_aic_0_targ_syscfg_apb_m_pready(i_aic_0_targ_syscfg_apb_m_pready),
        .o_aic_0_targ_syscfg_apb_m_psel(o_aic_0_targ_syscfg_apb_m_psel),
        .i_aic_0_targ_syscfg_apb_m_pslverr(i_aic_0_targ_syscfg_apb_m_pslverr),
        .o_aic_0_targ_syscfg_apb_m_pstrb(o_aic_0_targ_syscfg_apb_m_pstrb),
        .o_aic_0_targ_syscfg_apb_m_pwdata(o_aic_0_targ_syscfg_apb_m_pwdata),
        .o_aic_0_targ_syscfg_apb_m_pwrite(o_aic_0_targ_syscfg_apb_m_pwrite),
        .i_aic_1_aon_clk(i_aic_1_aon_clk),
        .i_aic_1_aon_rst_n(i_aic_1_aon_rst_n),
        .i_aic_1_clk(i_aic_1_clk),
        .i_aic_1_clken(i_aic_1_clken),
        .i_aic_1_init_ht_axi_s_araddr(i_aic_1_init_ht_axi_s_araddr),
        .i_aic_1_init_ht_axi_s_arburst(i_aic_1_init_ht_axi_s_arburst),
        .i_aic_1_init_ht_axi_s_arcache(i_aic_1_init_ht_axi_s_arcache),
        .i_aic_1_init_ht_axi_s_arid(i_aic_1_init_ht_axi_s_arid),
        .i_aic_1_init_ht_axi_s_arlen(i_aic_1_init_ht_axi_s_arlen),
        .i_aic_1_init_ht_axi_s_arlock(i_aic_1_init_ht_axi_s_arlock),
        .i_aic_1_init_ht_axi_s_arprot(i_aic_1_init_ht_axi_s_arprot),
        .o_aic_1_init_ht_axi_s_arready(o_aic_1_init_ht_axi_s_arready),
        .i_aic_1_init_ht_axi_s_arsize(i_aic_1_init_ht_axi_s_arsize),
        .i_aic_1_init_ht_axi_s_arvalid(i_aic_1_init_ht_axi_s_arvalid),
        .o_aic_1_init_ht_axi_s_rdata(o_aic_1_init_ht_axi_s_rdata),
        .o_aic_1_init_ht_axi_s_rid(o_aic_1_init_ht_axi_s_rid),
        .o_aic_1_init_ht_axi_s_rlast(o_aic_1_init_ht_axi_s_rlast),
        .i_aic_1_init_ht_axi_s_rready(i_aic_1_init_ht_axi_s_rready),
        .o_aic_1_init_ht_axi_s_rresp(o_aic_1_init_ht_axi_s_rresp),
        .o_aic_1_init_ht_axi_s_rvalid(o_aic_1_init_ht_axi_s_rvalid),
        .i_aic_1_init_ht_axi_s_awaddr(i_aic_1_init_ht_axi_s_awaddr),
        .i_aic_1_init_ht_axi_s_awburst(i_aic_1_init_ht_axi_s_awburst),
        .i_aic_1_init_ht_axi_s_awcache(i_aic_1_init_ht_axi_s_awcache),
        .i_aic_1_init_ht_axi_s_awid(i_aic_1_init_ht_axi_s_awid),
        .i_aic_1_init_ht_axi_s_awlen(i_aic_1_init_ht_axi_s_awlen),
        .i_aic_1_init_ht_axi_s_awlock(i_aic_1_init_ht_axi_s_awlock),
        .i_aic_1_init_ht_axi_s_awprot(i_aic_1_init_ht_axi_s_awprot),
        .o_aic_1_init_ht_axi_s_awready(o_aic_1_init_ht_axi_s_awready),
        .i_aic_1_init_ht_axi_s_awsize(i_aic_1_init_ht_axi_s_awsize),
        .i_aic_1_init_ht_axi_s_awvalid(i_aic_1_init_ht_axi_s_awvalid),
        .o_aic_1_init_ht_axi_s_bid(o_aic_1_init_ht_axi_s_bid),
        .i_aic_1_init_ht_axi_s_bready(i_aic_1_init_ht_axi_s_bready),
        .o_aic_1_init_ht_axi_s_bresp(o_aic_1_init_ht_axi_s_bresp),
        .o_aic_1_init_ht_axi_s_bvalid(o_aic_1_init_ht_axi_s_bvalid),
        .i_aic_1_init_ht_axi_s_wdata(i_aic_1_init_ht_axi_s_wdata),
        .i_aic_1_init_ht_axi_s_wlast(i_aic_1_init_ht_axi_s_wlast),
        .o_aic_1_init_ht_axi_s_wready(o_aic_1_init_ht_axi_s_wready),
        .i_aic_1_init_ht_axi_s_wstrb(i_aic_1_init_ht_axi_s_wstrb),
        .i_aic_1_init_ht_axi_s_wvalid(i_aic_1_init_ht_axi_s_wvalid),
        .i_aic_1_init_lt_axi_s_araddr(i_aic_1_init_lt_axi_s_araddr),
        .i_aic_1_init_lt_axi_s_arburst(i_aic_1_init_lt_axi_s_arburst),
        .i_aic_1_init_lt_axi_s_arcache(i_aic_1_init_lt_axi_s_arcache),
        .i_aic_1_init_lt_axi_s_arid(i_aic_1_init_lt_axi_s_arid),
        .i_aic_1_init_lt_axi_s_arlen(i_aic_1_init_lt_axi_s_arlen),
        .i_aic_1_init_lt_axi_s_arlock(i_aic_1_init_lt_axi_s_arlock),
        .i_aic_1_init_lt_axi_s_arprot(i_aic_1_init_lt_axi_s_arprot),
        .i_aic_1_init_lt_axi_s_arqos(i_aic_1_init_lt_axi_s_arqos),
        .o_aic_1_init_lt_axi_s_arready(o_aic_1_init_lt_axi_s_arready),
        .i_aic_1_init_lt_axi_s_arsize(i_aic_1_init_lt_axi_s_arsize),
        .i_aic_1_init_lt_axi_s_arvalid(i_aic_1_init_lt_axi_s_arvalid),
        .i_aic_1_init_lt_axi_s_awaddr(i_aic_1_init_lt_axi_s_awaddr),
        .i_aic_1_init_lt_axi_s_awburst(i_aic_1_init_lt_axi_s_awburst),
        .i_aic_1_init_lt_axi_s_awcache(i_aic_1_init_lt_axi_s_awcache),
        .i_aic_1_init_lt_axi_s_awid(i_aic_1_init_lt_axi_s_awid),
        .i_aic_1_init_lt_axi_s_awlen(i_aic_1_init_lt_axi_s_awlen),
        .i_aic_1_init_lt_axi_s_awlock(i_aic_1_init_lt_axi_s_awlock),
        .i_aic_1_init_lt_axi_s_awprot(i_aic_1_init_lt_axi_s_awprot),
        .i_aic_1_init_lt_axi_s_awqos(i_aic_1_init_lt_axi_s_awqos),
        .o_aic_1_init_lt_axi_s_awready(o_aic_1_init_lt_axi_s_awready),
        .i_aic_1_init_lt_axi_s_awsize(i_aic_1_init_lt_axi_s_awsize),
        .i_aic_1_init_lt_axi_s_awvalid(i_aic_1_init_lt_axi_s_awvalid),
        .o_aic_1_init_lt_axi_s_bid(o_aic_1_init_lt_axi_s_bid),
        .i_aic_1_init_lt_axi_s_bready(i_aic_1_init_lt_axi_s_bready),
        .o_aic_1_init_lt_axi_s_bresp(o_aic_1_init_lt_axi_s_bresp),
        .o_aic_1_init_lt_axi_s_bvalid(o_aic_1_init_lt_axi_s_bvalid),
        .o_aic_1_init_lt_axi_s_rdata(o_aic_1_init_lt_axi_s_rdata),
        .o_aic_1_init_lt_axi_s_rid(o_aic_1_init_lt_axi_s_rid),
        .o_aic_1_init_lt_axi_s_rlast(o_aic_1_init_lt_axi_s_rlast),
        .i_aic_1_init_lt_axi_s_rready(i_aic_1_init_lt_axi_s_rready),
        .o_aic_1_init_lt_axi_s_rresp(o_aic_1_init_lt_axi_s_rresp),
        .o_aic_1_init_lt_axi_s_rvalid(o_aic_1_init_lt_axi_s_rvalid),
        .i_aic_1_init_lt_axi_s_wdata(i_aic_1_init_lt_axi_s_wdata),
        .i_aic_1_init_lt_axi_s_wlast(i_aic_1_init_lt_axi_s_wlast),
        .o_aic_1_init_lt_axi_s_wready(o_aic_1_init_lt_axi_s_wready),
        .i_aic_1_init_lt_axi_s_wstrb(i_aic_1_init_lt_axi_s_wstrb),
        .i_aic_1_init_lt_axi_s_wvalid(i_aic_1_init_lt_axi_s_wvalid),
        .o_aic_1_pwr_idle_val(o_aic_1_pwr_idle_val),
        .o_aic_1_pwr_idle_ack(o_aic_1_pwr_idle_ack),
        .i_aic_1_pwr_idle_req(i_aic_1_pwr_idle_req),
        .i_aic_1_rst_n(i_aic_1_rst_n),
        .o_aic_1_targ_lt_axi_m_araddr(o_aic_1_targ_lt_axi_m_araddr),
        .o_aic_1_targ_lt_axi_m_arburst(o_aic_1_targ_lt_axi_m_arburst),
        .o_aic_1_targ_lt_axi_m_arcache(o_aic_1_targ_lt_axi_m_arcache),
        .o_aic_1_targ_lt_axi_m_arid(o_aic_1_targ_lt_axi_m_arid),
        .o_aic_1_targ_lt_axi_m_arlen(o_aic_1_targ_lt_axi_m_arlen),
        .o_aic_1_targ_lt_axi_m_arlock(o_aic_1_targ_lt_axi_m_arlock),
        .o_aic_1_targ_lt_axi_m_arprot(o_aic_1_targ_lt_axi_m_arprot),
        .o_aic_1_targ_lt_axi_m_arqos(o_aic_1_targ_lt_axi_m_arqos),
        .i_aic_1_targ_lt_axi_m_arready(i_aic_1_targ_lt_axi_m_arready),
        .o_aic_1_targ_lt_axi_m_arsize(o_aic_1_targ_lt_axi_m_arsize),
        .o_aic_1_targ_lt_axi_m_arvalid(o_aic_1_targ_lt_axi_m_arvalid),
        .o_aic_1_targ_lt_axi_m_awaddr(o_aic_1_targ_lt_axi_m_awaddr),
        .o_aic_1_targ_lt_axi_m_awburst(o_aic_1_targ_lt_axi_m_awburst),
        .o_aic_1_targ_lt_axi_m_awcache(o_aic_1_targ_lt_axi_m_awcache),
        .o_aic_1_targ_lt_axi_m_awid(o_aic_1_targ_lt_axi_m_awid),
        .o_aic_1_targ_lt_axi_m_awlen(o_aic_1_targ_lt_axi_m_awlen),
        .o_aic_1_targ_lt_axi_m_awlock(o_aic_1_targ_lt_axi_m_awlock),
        .o_aic_1_targ_lt_axi_m_awprot(o_aic_1_targ_lt_axi_m_awprot),
        .o_aic_1_targ_lt_axi_m_awqos(o_aic_1_targ_lt_axi_m_awqos),
        .i_aic_1_targ_lt_axi_m_awready(i_aic_1_targ_lt_axi_m_awready),
        .o_aic_1_targ_lt_axi_m_awsize(o_aic_1_targ_lt_axi_m_awsize),
        .o_aic_1_targ_lt_axi_m_awvalid(o_aic_1_targ_lt_axi_m_awvalid),
        .i_aic_1_targ_lt_axi_m_bid(i_aic_1_targ_lt_axi_m_bid),
        .o_aic_1_targ_lt_axi_m_bready(o_aic_1_targ_lt_axi_m_bready),
        .i_aic_1_targ_lt_axi_m_bresp(i_aic_1_targ_lt_axi_m_bresp),
        .i_aic_1_targ_lt_axi_m_bvalid(i_aic_1_targ_lt_axi_m_bvalid),
        .i_aic_1_targ_lt_axi_m_rdata(i_aic_1_targ_lt_axi_m_rdata),
        .i_aic_1_targ_lt_axi_m_rid(i_aic_1_targ_lt_axi_m_rid),
        .i_aic_1_targ_lt_axi_m_rlast(i_aic_1_targ_lt_axi_m_rlast),
        .o_aic_1_targ_lt_axi_m_rready(o_aic_1_targ_lt_axi_m_rready),
        .i_aic_1_targ_lt_axi_m_rresp(i_aic_1_targ_lt_axi_m_rresp),
        .i_aic_1_targ_lt_axi_m_rvalid(i_aic_1_targ_lt_axi_m_rvalid),
        .o_aic_1_targ_lt_axi_m_wdata(o_aic_1_targ_lt_axi_m_wdata),
        .o_aic_1_targ_lt_axi_m_wlast(o_aic_1_targ_lt_axi_m_wlast),
        .i_aic_1_targ_lt_axi_m_wready(i_aic_1_targ_lt_axi_m_wready),
        .o_aic_1_targ_lt_axi_m_wstrb(o_aic_1_targ_lt_axi_m_wstrb),
        .o_aic_1_targ_lt_axi_m_wvalid(o_aic_1_targ_lt_axi_m_wvalid),
        .o_aic_1_targ_syscfg_apb_m_paddr(o_aic_1_targ_syscfg_apb_m_paddr),
        .o_aic_1_targ_syscfg_apb_m_penable(o_aic_1_targ_syscfg_apb_m_penable),
        .o_aic_1_targ_syscfg_apb_m_pprot(o_aic_1_targ_syscfg_apb_m_pprot),
        .i_aic_1_targ_syscfg_apb_m_prdata(i_aic_1_targ_syscfg_apb_m_prdata),
        .i_aic_1_targ_syscfg_apb_m_pready(i_aic_1_targ_syscfg_apb_m_pready),
        .o_aic_1_targ_syscfg_apb_m_psel(o_aic_1_targ_syscfg_apb_m_psel),
        .i_aic_1_targ_syscfg_apb_m_pslverr(i_aic_1_targ_syscfg_apb_m_pslverr),
        .o_aic_1_targ_syscfg_apb_m_pstrb(o_aic_1_targ_syscfg_apb_m_pstrb),
        .o_aic_1_targ_syscfg_apb_m_pwdata(o_aic_1_targ_syscfg_apb_m_pwdata),
        .o_aic_1_targ_syscfg_apb_m_pwrite(o_aic_1_targ_syscfg_apb_m_pwrite),
        .i_aic_2_aon_clk(i_aic_2_aon_clk),
        .i_aic_2_aon_rst_n(i_aic_2_aon_rst_n),
        .i_aic_2_clk(i_aic_2_clk),
        .i_aic_2_clken(i_aic_2_clken),
        .i_aic_2_init_ht_axi_s_araddr(i_aic_2_init_ht_axi_s_araddr),
        .i_aic_2_init_ht_axi_s_arburst(i_aic_2_init_ht_axi_s_arburst),
        .i_aic_2_init_ht_axi_s_arcache(i_aic_2_init_ht_axi_s_arcache),
        .i_aic_2_init_ht_axi_s_arid(i_aic_2_init_ht_axi_s_arid),
        .i_aic_2_init_ht_axi_s_arlen(i_aic_2_init_ht_axi_s_arlen),
        .i_aic_2_init_ht_axi_s_arlock(i_aic_2_init_ht_axi_s_arlock),
        .i_aic_2_init_ht_axi_s_arprot(i_aic_2_init_ht_axi_s_arprot),
        .o_aic_2_init_ht_axi_s_arready(o_aic_2_init_ht_axi_s_arready),
        .i_aic_2_init_ht_axi_s_arsize(i_aic_2_init_ht_axi_s_arsize),
        .i_aic_2_init_ht_axi_s_arvalid(i_aic_2_init_ht_axi_s_arvalid),
        .o_aic_2_init_ht_axi_s_rdata(o_aic_2_init_ht_axi_s_rdata),
        .o_aic_2_init_ht_axi_s_rid(o_aic_2_init_ht_axi_s_rid),
        .o_aic_2_init_ht_axi_s_rlast(o_aic_2_init_ht_axi_s_rlast),
        .i_aic_2_init_ht_axi_s_rready(i_aic_2_init_ht_axi_s_rready),
        .o_aic_2_init_ht_axi_s_rresp(o_aic_2_init_ht_axi_s_rresp),
        .o_aic_2_init_ht_axi_s_rvalid(o_aic_2_init_ht_axi_s_rvalid),
        .i_aic_2_init_ht_axi_s_awaddr(i_aic_2_init_ht_axi_s_awaddr),
        .i_aic_2_init_ht_axi_s_awburst(i_aic_2_init_ht_axi_s_awburst),
        .i_aic_2_init_ht_axi_s_awcache(i_aic_2_init_ht_axi_s_awcache),
        .i_aic_2_init_ht_axi_s_awid(i_aic_2_init_ht_axi_s_awid),
        .i_aic_2_init_ht_axi_s_awlen(i_aic_2_init_ht_axi_s_awlen),
        .i_aic_2_init_ht_axi_s_awlock(i_aic_2_init_ht_axi_s_awlock),
        .i_aic_2_init_ht_axi_s_awprot(i_aic_2_init_ht_axi_s_awprot),
        .o_aic_2_init_ht_axi_s_awready(o_aic_2_init_ht_axi_s_awready),
        .i_aic_2_init_ht_axi_s_awsize(i_aic_2_init_ht_axi_s_awsize),
        .i_aic_2_init_ht_axi_s_awvalid(i_aic_2_init_ht_axi_s_awvalid),
        .o_aic_2_init_ht_axi_s_bid(o_aic_2_init_ht_axi_s_bid),
        .i_aic_2_init_ht_axi_s_bready(i_aic_2_init_ht_axi_s_bready),
        .o_aic_2_init_ht_axi_s_bresp(o_aic_2_init_ht_axi_s_bresp),
        .o_aic_2_init_ht_axi_s_bvalid(o_aic_2_init_ht_axi_s_bvalid),
        .i_aic_2_init_ht_axi_s_wdata(i_aic_2_init_ht_axi_s_wdata),
        .i_aic_2_init_ht_axi_s_wlast(i_aic_2_init_ht_axi_s_wlast),
        .o_aic_2_init_ht_axi_s_wready(o_aic_2_init_ht_axi_s_wready),
        .i_aic_2_init_ht_axi_s_wstrb(i_aic_2_init_ht_axi_s_wstrb),
        .i_aic_2_init_ht_axi_s_wvalid(i_aic_2_init_ht_axi_s_wvalid),
        .i_aic_2_init_lt_axi_s_araddr(i_aic_2_init_lt_axi_s_araddr),
        .i_aic_2_init_lt_axi_s_arburst(i_aic_2_init_lt_axi_s_arburst),
        .i_aic_2_init_lt_axi_s_arcache(i_aic_2_init_lt_axi_s_arcache),
        .i_aic_2_init_lt_axi_s_arid(i_aic_2_init_lt_axi_s_arid),
        .i_aic_2_init_lt_axi_s_arlen(i_aic_2_init_lt_axi_s_arlen),
        .i_aic_2_init_lt_axi_s_arlock(i_aic_2_init_lt_axi_s_arlock),
        .i_aic_2_init_lt_axi_s_arprot(i_aic_2_init_lt_axi_s_arprot),
        .i_aic_2_init_lt_axi_s_arqos(i_aic_2_init_lt_axi_s_arqos),
        .o_aic_2_init_lt_axi_s_arready(o_aic_2_init_lt_axi_s_arready),
        .i_aic_2_init_lt_axi_s_arsize(i_aic_2_init_lt_axi_s_arsize),
        .i_aic_2_init_lt_axi_s_arvalid(i_aic_2_init_lt_axi_s_arvalid),
        .i_aic_2_init_lt_axi_s_awaddr(i_aic_2_init_lt_axi_s_awaddr),
        .i_aic_2_init_lt_axi_s_awburst(i_aic_2_init_lt_axi_s_awburst),
        .i_aic_2_init_lt_axi_s_awcache(i_aic_2_init_lt_axi_s_awcache),
        .i_aic_2_init_lt_axi_s_awid(i_aic_2_init_lt_axi_s_awid),
        .i_aic_2_init_lt_axi_s_awlen(i_aic_2_init_lt_axi_s_awlen),
        .i_aic_2_init_lt_axi_s_awlock(i_aic_2_init_lt_axi_s_awlock),
        .i_aic_2_init_lt_axi_s_awprot(i_aic_2_init_lt_axi_s_awprot),
        .i_aic_2_init_lt_axi_s_awqos(i_aic_2_init_lt_axi_s_awqos),
        .o_aic_2_init_lt_axi_s_awready(o_aic_2_init_lt_axi_s_awready),
        .i_aic_2_init_lt_axi_s_awsize(i_aic_2_init_lt_axi_s_awsize),
        .i_aic_2_init_lt_axi_s_awvalid(i_aic_2_init_lt_axi_s_awvalid),
        .o_aic_2_init_lt_axi_s_bid(o_aic_2_init_lt_axi_s_bid),
        .i_aic_2_init_lt_axi_s_bready(i_aic_2_init_lt_axi_s_bready),
        .o_aic_2_init_lt_axi_s_bresp(o_aic_2_init_lt_axi_s_bresp),
        .o_aic_2_init_lt_axi_s_bvalid(o_aic_2_init_lt_axi_s_bvalid),
        .o_aic_2_init_lt_axi_s_rdata(o_aic_2_init_lt_axi_s_rdata),
        .o_aic_2_init_lt_axi_s_rid(o_aic_2_init_lt_axi_s_rid),
        .o_aic_2_init_lt_axi_s_rlast(o_aic_2_init_lt_axi_s_rlast),
        .i_aic_2_init_lt_axi_s_rready(i_aic_2_init_lt_axi_s_rready),
        .o_aic_2_init_lt_axi_s_rresp(o_aic_2_init_lt_axi_s_rresp),
        .o_aic_2_init_lt_axi_s_rvalid(o_aic_2_init_lt_axi_s_rvalid),
        .i_aic_2_init_lt_axi_s_wdata(i_aic_2_init_lt_axi_s_wdata),
        .i_aic_2_init_lt_axi_s_wlast(i_aic_2_init_lt_axi_s_wlast),
        .o_aic_2_init_lt_axi_s_wready(o_aic_2_init_lt_axi_s_wready),
        .i_aic_2_init_lt_axi_s_wstrb(i_aic_2_init_lt_axi_s_wstrb),
        .i_aic_2_init_lt_axi_s_wvalid(i_aic_2_init_lt_axi_s_wvalid),
        .o_aic_2_pwr_idle_val(o_aic_2_pwr_idle_val),
        .o_aic_2_pwr_idle_ack(o_aic_2_pwr_idle_ack),
        .i_aic_2_pwr_idle_req(i_aic_2_pwr_idle_req),
        .i_aic_2_rst_n(i_aic_2_rst_n),
        .o_aic_2_targ_lt_axi_m_araddr(o_aic_2_targ_lt_axi_m_araddr),
        .o_aic_2_targ_lt_axi_m_arburst(o_aic_2_targ_lt_axi_m_arburst),
        .o_aic_2_targ_lt_axi_m_arcache(o_aic_2_targ_lt_axi_m_arcache),
        .o_aic_2_targ_lt_axi_m_arid(o_aic_2_targ_lt_axi_m_arid),
        .o_aic_2_targ_lt_axi_m_arlen(o_aic_2_targ_lt_axi_m_arlen),
        .o_aic_2_targ_lt_axi_m_arlock(o_aic_2_targ_lt_axi_m_arlock),
        .o_aic_2_targ_lt_axi_m_arprot(o_aic_2_targ_lt_axi_m_arprot),
        .o_aic_2_targ_lt_axi_m_arqos(o_aic_2_targ_lt_axi_m_arqos),
        .i_aic_2_targ_lt_axi_m_arready(i_aic_2_targ_lt_axi_m_arready),
        .o_aic_2_targ_lt_axi_m_arsize(o_aic_2_targ_lt_axi_m_arsize),
        .o_aic_2_targ_lt_axi_m_arvalid(o_aic_2_targ_lt_axi_m_arvalid),
        .o_aic_2_targ_lt_axi_m_awaddr(o_aic_2_targ_lt_axi_m_awaddr),
        .o_aic_2_targ_lt_axi_m_awburst(o_aic_2_targ_lt_axi_m_awburst),
        .o_aic_2_targ_lt_axi_m_awcache(o_aic_2_targ_lt_axi_m_awcache),
        .o_aic_2_targ_lt_axi_m_awid(o_aic_2_targ_lt_axi_m_awid),
        .o_aic_2_targ_lt_axi_m_awlen(o_aic_2_targ_lt_axi_m_awlen),
        .o_aic_2_targ_lt_axi_m_awlock(o_aic_2_targ_lt_axi_m_awlock),
        .o_aic_2_targ_lt_axi_m_awprot(o_aic_2_targ_lt_axi_m_awprot),
        .o_aic_2_targ_lt_axi_m_awqos(o_aic_2_targ_lt_axi_m_awqos),
        .i_aic_2_targ_lt_axi_m_awready(i_aic_2_targ_lt_axi_m_awready),
        .o_aic_2_targ_lt_axi_m_awsize(o_aic_2_targ_lt_axi_m_awsize),
        .o_aic_2_targ_lt_axi_m_awvalid(o_aic_2_targ_lt_axi_m_awvalid),
        .i_aic_2_targ_lt_axi_m_bid(i_aic_2_targ_lt_axi_m_bid),
        .o_aic_2_targ_lt_axi_m_bready(o_aic_2_targ_lt_axi_m_bready),
        .i_aic_2_targ_lt_axi_m_bresp(i_aic_2_targ_lt_axi_m_bresp),
        .i_aic_2_targ_lt_axi_m_bvalid(i_aic_2_targ_lt_axi_m_bvalid),
        .i_aic_2_targ_lt_axi_m_rdata(i_aic_2_targ_lt_axi_m_rdata),
        .i_aic_2_targ_lt_axi_m_rid(i_aic_2_targ_lt_axi_m_rid),
        .i_aic_2_targ_lt_axi_m_rlast(i_aic_2_targ_lt_axi_m_rlast),
        .o_aic_2_targ_lt_axi_m_rready(o_aic_2_targ_lt_axi_m_rready),
        .i_aic_2_targ_lt_axi_m_rresp(i_aic_2_targ_lt_axi_m_rresp),
        .i_aic_2_targ_lt_axi_m_rvalid(i_aic_2_targ_lt_axi_m_rvalid),
        .o_aic_2_targ_lt_axi_m_wdata(o_aic_2_targ_lt_axi_m_wdata),
        .o_aic_2_targ_lt_axi_m_wlast(o_aic_2_targ_lt_axi_m_wlast),
        .i_aic_2_targ_lt_axi_m_wready(i_aic_2_targ_lt_axi_m_wready),
        .o_aic_2_targ_lt_axi_m_wstrb(o_aic_2_targ_lt_axi_m_wstrb),
        .o_aic_2_targ_lt_axi_m_wvalid(o_aic_2_targ_lt_axi_m_wvalid),
        .o_aic_2_targ_syscfg_apb_m_paddr(o_aic_2_targ_syscfg_apb_m_paddr),
        .o_aic_2_targ_syscfg_apb_m_penable(o_aic_2_targ_syscfg_apb_m_penable),
        .o_aic_2_targ_syscfg_apb_m_pprot(o_aic_2_targ_syscfg_apb_m_pprot),
        .i_aic_2_targ_syscfg_apb_m_prdata(i_aic_2_targ_syscfg_apb_m_prdata),
        .i_aic_2_targ_syscfg_apb_m_pready(i_aic_2_targ_syscfg_apb_m_pready),
        .o_aic_2_targ_syscfg_apb_m_psel(o_aic_2_targ_syscfg_apb_m_psel),
        .i_aic_2_targ_syscfg_apb_m_pslverr(i_aic_2_targ_syscfg_apb_m_pslverr),
        .o_aic_2_targ_syscfg_apb_m_pstrb(o_aic_2_targ_syscfg_apb_m_pstrb),
        .o_aic_2_targ_syscfg_apb_m_pwdata(o_aic_2_targ_syscfg_apb_m_pwdata),
        .o_aic_2_targ_syscfg_apb_m_pwrite(o_aic_2_targ_syscfg_apb_m_pwrite),
        .i_aic_3_aon_clk(i_aic_3_aon_clk),
        .i_aic_3_aon_rst_n(i_aic_3_aon_rst_n),
        .i_aic_3_clk(i_aic_3_clk),
        .i_aic_3_clken(i_aic_3_clken),
        .i_aic_3_init_ht_axi_s_araddr(i_aic_3_init_ht_axi_s_araddr),
        .i_aic_3_init_ht_axi_s_arburst(i_aic_3_init_ht_axi_s_arburst),
        .i_aic_3_init_ht_axi_s_arcache(i_aic_3_init_ht_axi_s_arcache),
        .i_aic_3_init_ht_axi_s_arid(i_aic_3_init_ht_axi_s_arid),
        .i_aic_3_init_ht_axi_s_arlen(i_aic_3_init_ht_axi_s_arlen),
        .i_aic_3_init_ht_axi_s_arlock(i_aic_3_init_ht_axi_s_arlock),
        .i_aic_3_init_ht_axi_s_arprot(i_aic_3_init_ht_axi_s_arprot),
        .o_aic_3_init_ht_axi_s_arready(o_aic_3_init_ht_axi_s_arready),
        .i_aic_3_init_ht_axi_s_arsize(i_aic_3_init_ht_axi_s_arsize),
        .i_aic_3_init_ht_axi_s_arvalid(i_aic_3_init_ht_axi_s_arvalid),
        .o_aic_3_init_ht_axi_s_rdata(o_aic_3_init_ht_axi_s_rdata),
        .o_aic_3_init_ht_axi_s_rid(o_aic_3_init_ht_axi_s_rid),
        .o_aic_3_init_ht_axi_s_rlast(o_aic_3_init_ht_axi_s_rlast),
        .i_aic_3_init_ht_axi_s_rready(i_aic_3_init_ht_axi_s_rready),
        .o_aic_3_init_ht_axi_s_rresp(o_aic_3_init_ht_axi_s_rresp),
        .o_aic_3_init_ht_axi_s_rvalid(o_aic_3_init_ht_axi_s_rvalid),
        .i_aic_3_init_ht_axi_s_awaddr(i_aic_3_init_ht_axi_s_awaddr),
        .i_aic_3_init_ht_axi_s_awburst(i_aic_3_init_ht_axi_s_awburst),
        .i_aic_3_init_ht_axi_s_awcache(i_aic_3_init_ht_axi_s_awcache),
        .i_aic_3_init_ht_axi_s_awid(i_aic_3_init_ht_axi_s_awid),
        .i_aic_3_init_ht_axi_s_awlen(i_aic_3_init_ht_axi_s_awlen),
        .i_aic_3_init_ht_axi_s_awlock(i_aic_3_init_ht_axi_s_awlock),
        .i_aic_3_init_ht_axi_s_awprot(i_aic_3_init_ht_axi_s_awprot),
        .o_aic_3_init_ht_axi_s_awready(o_aic_3_init_ht_axi_s_awready),
        .i_aic_3_init_ht_axi_s_awsize(i_aic_3_init_ht_axi_s_awsize),
        .i_aic_3_init_ht_axi_s_awvalid(i_aic_3_init_ht_axi_s_awvalid),
        .o_aic_3_init_ht_axi_s_bid(o_aic_3_init_ht_axi_s_bid),
        .i_aic_3_init_ht_axi_s_bready(i_aic_3_init_ht_axi_s_bready),
        .o_aic_3_init_ht_axi_s_bresp(o_aic_3_init_ht_axi_s_bresp),
        .o_aic_3_init_ht_axi_s_bvalid(o_aic_3_init_ht_axi_s_bvalid),
        .i_aic_3_init_ht_axi_s_wdata(i_aic_3_init_ht_axi_s_wdata),
        .i_aic_3_init_ht_axi_s_wlast(i_aic_3_init_ht_axi_s_wlast),
        .o_aic_3_init_ht_axi_s_wready(o_aic_3_init_ht_axi_s_wready),
        .i_aic_3_init_ht_axi_s_wstrb(i_aic_3_init_ht_axi_s_wstrb),
        .i_aic_3_init_ht_axi_s_wvalid(i_aic_3_init_ht_axi_s_wvalid),
        .i_aic_3_init_lt_axi_s_araddr(i_aic_3_init_lt_axi_s_araddr),
        .i_aic_3_init_lt_axi_s_arburst(i_aic_3_init_lt_axi_s_arburst),
        .i_aic_3_init_lt_axi_s_arcache(i_aic_3_init_lt_axi_s_arcache),
        .i_aic_3_init_lt_axi_s_arid(i_aic_3_init_lt_axi_s_arid),
        .i_aic_3_init_lt_axi_s_arlen(i_aic_3_init_lt_axi_s_arlen),
        .i_aic_3_init_lt_axi_s_arlock(i_aic_3_init_lt_axi_s_arlock),
        .i_aic_3_init_lt_axi_s_arprot(i_aic_3_init_lt_axi_s_arprot),
        .i_aic_3_init_lt_axi_s_arqos(i_aic_3_init_lt_axi_s_arqos),
        .o_aic_3_init_lt_axi_s_arready(o_aic_3_init_lt_axi_s_arready),
        .i_aic_3_init_lt_axi_s_arsize(i_aic_3_init_lt_axi_s_arsize),
        .i_aic_3_init_lt_axi_s_arvalid(i_aic_3_init_lt_axi_s_arvalid),
        .i_aic_3_init_lt_axi_s_awaddr(i_aic_3_init_lt_axi_s_awaddr),
        .i_aic_3_init_lt_axi_s_awburst(i_aic_3_init_lt_axi_s_awburst),
        .i_aic_3_init_lt_axi_s_awcache(i_aic_3_init_lt_axi_s_awcache),
        .i_aic_3_init_lt_axi_s_awid(i_aic_3_init_lt_axi_s_awid),
        .i_aic_3_init_lt_axi_s_awlen(i_aic_3_init_lt_axi_s_awlen),
        .i_aic_3_init_lt_axi_s_awlock(i_aic_3_init_lt_axi_s_awlock),
        .i_aic_3_init_lt_axi_s_awprot(i_aic_3_init_lt_axi_s_awprot),
        .i_aic_3_init_lt_axi_s_awqos(i_aic_3_init_lt_axi_s_awqos),
        .o_aic_3_init_lt_axi_s_awready(o_aic_3_init_lt_axi_s_awready),
        .i_aic_3_init_lt_axi_s_awsize(i_aic_3_init_lt_axi_s_awsize),
        .i_aic_3_init_lt_axi_s_awvalid(i_aic_3_init_lt_axi_s_awvalid),
        .o_aic_3_init_lt_axi_s_bid(o_aic_3_init_lt_axi_s_bid),
        .i_aic_3_init_lt_axi_s_bready(i_aic_3_init_lt_axi_s_bready),
        .o_aic_3_init_lt_axi_s_bresp(o_aic_3_init_lt_axi_s_bresp),
        .o_aic_3_init_lt_axi_s_bvalid(o_aic_3_init_lt_axi_s_bvalid),
        .o_aic_3_init_lt_axi_s_rdata(o_aic_3_init_lt_axi_s_rdata),
        .o_aic_3_init_lt_axi_s_rid(o_aic_3_init_lt_axi_s_rid),
        .o_aic_3_init_lt_axi_s_rlast(o_aic_3_init_lt_axi_s_rlast),
        .i_aic_3_init_lt_axi_s_rready(i_aic_3_init_lt_axi_s_rready),
        .o_aic_3_init_lt_axi_s_rresp(o_aic_3_init_lt_axi_s_rresp),
        .o_aic_3_init_lt_axi_s_rvalid(o_aic_3_init_lt_axi_s_rvalid),
        .i_aic_3_init_lt_axi_s_wdata(i_aic_3_init_lt_axi_s_wdata),
        .i_aic_3_init_lt_axi_s_wlast(i_aic_3_init_lt_axi_s_wlast),
        .o_aic_3_init_lt_axi_s_wready(o_aic_3_init_lt_axi_s_wready),
        .i_aic_3_init_lt_axi_s_wstrb(i_aic_3_init_lt_axi_s_wstrb),
        .i_aic_3_init_lt_axi_s_wvalid(i_aic_3_init_lt_axi_s_wvalid),
        .i_aic_3_init_tok_ocpl_s_maddr(i_aic_3_init_tok_ocpl_s_maddr),
        .i_aic_3_init_tok_ocpl_s_mcmd(i_aic_3_init_tok_ocpl_s_mcmd),
        .i_aic_3_init_tok_ocpl_s_mdata(i_aic_3_init_tok_ocpl_s_mdata),
        .o_aic_3_init_tok_ocpl_s_scmdaccept(o_aic_3_init_tok_ocpl_s_scmdaccept),
        .o_aic_3_pwr_idle_val(o_aic_3_pwr_idle_val),
        .o_aic_3_pwr_idle_ack(o_aic_3_pwr_idle_ack),
        .i_aic_3_pwr_idle_req(i_aic_3_pwr_idle_req),
        .i_aic_3_rst_n(i_aic_3_rst_n),
        .o_aic_3_targ_lt_axi_m_araddr(o_aic_3_targ_lt_axi_m_araddr),
        .o_aic_3_targ_lt_axi_m_arburst(o_aic_3_targ_lt_axi_m_arburst),
        .o_aic_3_targ_lt_axi_m_arcache(o_aic_3_targ_lt_axi_m_arcache),
        .o_aic_3_targ_lt_axi_m_arid(o_aic_3_targ_lt_axi_m_arid),
        .o_aic_3_targ_lt_axi_m_arlen(o_aic_3_targ_lt_axi_m_arlen),
        .o_aic_3_targ_lt_axi_m_arlock(o_aic_3_targ_lt_axi_m_arlock),
        .o_aic_3_targ_lt_axi_m_arprot(o_aic_3_targ_lt_axi_m_arprot),
        .o_aic_3_targ_lt_axi_m_arqos(o_aic_3_targ_lt_axi_m_arqos),
        .i_aic_3_targ_lt_axi_m_arready(i_aic_3_targ_lt_axi_m_arready),
        .o_aic_3_targ_lt_axi_m_arsize(o_aic_3_targ_lt_axi_m_arsize),
        .o_aic_3_targ_lt_axi_m_arvalid(o_aic_3_targ_lt_axi_m_arvalid),
        .o_aic_3_targ_lt_axi_m_awaddr(o_aic_3_targ_lt_axi_m_awaddr),
        .o_aic_3_targ_lt_axi_m_awburst(o_aic_3_targ_lt_axi_m_awburst),
        .o_aic_3_targ_lt_axi_m_awcache(o_aic_3_targ_lt_axi_m_awcache),
        .o_aic_3_targ_lt_axi_m_awid(o_aic_3_targ_lt_axi_m_awid),
        .o_aic_3_targ_lt_axi_m_awlen(o_aic_3_targ_lt_axi_m_awlen),
        .o_aic_3_targ_lt_axi_m_awlock(o_aic_3_targ_lt_axi_m_awlock),
        .o_aic_3_targ_lt_axi_m_awprot(o_aic_3_targ_lt_axi_m_awprot),
        .o_aic_3_targ_lt_axi_m_awqos(o_aic_3_targ_lt_axi_m_awqos),
        .i_aic_3_targ_lt_axi_m_awready(i_aic_3_targ_lt_axi_m_awready),
        .o_aic_3_targ_lt_axi_m_awsize(o_aic_3_targ_lt_axi_m_awsize),
        .o_aic_3_targ_lt_axi_m_awvalid(o_aic_3_targ_lt_axi_m_awvalid),
        .i_aic_3_targ_lt_axi_m_bid(i_aic_3_targ_lt_axi_m_bid),
        .o_aic_3_targ_lt_axi_m_bready(o_aic_3_targ_lt_axi_m_bready),
        .i_aic_3_targ_lt_axi_m_bresp(i_aic_3_targ_lt_axi_m_bresp),
        .i_aic_3_targ_lt_axi_m_bvalid(i_aic_3_targ_lt_axi_m_bvalid),
        .i_aic_3_targ_lt_axi_m_rdata(i_aic_3_targ_lt_axi_m_rdata),
        .i_aic_3_targ_lt_axi_m_rid(i_aic_3_targ_lt_axi_m_rid),
        .i_aic_3_targ_lt_axi_m_rlast(i_aic_3_targ_lt_axi_m_rlast),
        .o_aic_3_targ_lt_axi_m_rready(o_aic_3_targ_lt_axi_m_rready),
        .i_aic_3_targ_lt_axi_m_rresp(i_aic_3_targ_lt_axi_m_rresp),
        .i_aic_3_targ_lt_axi_m_rvalid(i_aic_3_targ_lt_axi_m_rvalid),
        .o_aic_3_targ_lt_axi_m_wdata(o_aic_3_targ_lt_axi_m_wdata),
        .o_aic_3_targ_lt_axi_m_wlast(o_aic_3_targ_lt_axi_m_wlast),
        .i_aic_3_targ_lt_axi_m_wready(i_aic_3_targ_lt_axi_m_wready),
        .o_aic_3_targ_lt_axi_m_wstrb(o_aic_3_targ_lt_axi_m_wstrb),
        .o_aic_3_targ_lt_axi_m_wvalid(o_aic_3_targ_lt_axi_m_wvalid),
        .o_aic_3_targ_syscfg_apb_m_paddr(o_aic_3_targ_syscfg_apb_m_paddr),
        .o_aic_3_targ_syscfg_apb_m_penable(o_aic_3_targ_syscfg_apb_m_penable),
        .o_aic_3_targ_syscfg_apb_m_pprot(o_aic_3_targ_syscfg_apb_m_pprot),
        .i_aic_3_targ_syscfg_apb_m_prdata(i_aic_3_targ_syscfg_apb_m_prdata),
        .i_aic_3_targ_syscfg_apb_m_pready(i_aic_3_targ_syscfg_apb_m_pready),
        .o_aic_3_targ_syscfg_apb_m_psel(o_aic_3_targ_syscfg_apb_m_psel),
        .i_aic_3_targ_syscfg_apb_m_pslverr(i_aic_3_targ_syscfg_apb_m_pslverr),
        .o_aic_3_targ_syscfg_apb_m_pstrb(o_aic_3_targ_syscfg_apb_m_pstrb),
        .o_aic_3_targ_syscfg_apb_m_pwdata(o_aic_3_targ_syscfg_apb_m_pwdata),
        .o_aic_3_targ_syscfg_apb_m_pwrite(o_aic_3_targ_syscfg_apb_m_pwrite),
        .i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data),
        .i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head),
        .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail),
        .i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld),
        .o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data),
        .i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head),
        .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy),
        .i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail),
        .i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld),
        .o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data),
        .o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head),
        .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data),
        .i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head),
        .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy),
        .i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail),
        .i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld),
        .o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data),
        .o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head),
        .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail),
        .o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data),
        .o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head),
        .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail),
        .o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld),
        .i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data),
        .o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head),
        .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail),
        .o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld),
        .i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data),
        .o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head),
        .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail),
        .o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld),
        .i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data),
        .o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head),
        .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail),
        .o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld),
        .i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data),
        .o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head),
        .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail),
        .o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld),
        .i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data),
        .o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head),
        .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail),
        .o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld),
        .i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data),
        .o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head),
        .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail),
        .o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld),
        .i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data),
        .o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head),
        .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail),
        .o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld),
        .i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data),
        .o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head),
        .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail),
        .o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld),
        .i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data),
        .o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head),
        .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail),
        .o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld),
        .i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data),
        .o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head),
        .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail),
        .o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld),
        .i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data),
        .o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head),
        .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy),
        .o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail),
        .o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld),
        .i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data),
        .i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head),
        .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data),
        .o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head),
        .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy),
        .o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail),
        .o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld),
        .i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data),
        .i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head),
        .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail),
        .i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld),
        .i_l2_0_aon_clk(i_l2_0_aon_clk),
        .i_l2_0_aon_rst_n(i_l2_0_aon_rst_n),
        .i_l2_0_clk(i_l2_0_clk),
        .i_l2_0_clken(i_l2_0_clken),
        .o_l2_0_pwr_idle_val(o_l2_0_pwr_idle_val),
        .o_l2_0_pwr_idle_ack(o_l2_0_pwr_idle_ack),
        .i_l2_0_pwr_idle_req(i_l2_0_pwr_idle_req),
        .i_l2_0_rst_n(i_l2_0_rst_n),
        .o_l2_0_targ_ht_axi_m_araddr(o_l2_0_targ_ht_axi_m_araddr),
        .o_l2_0_targ_ht_axi_m_arburst(o_l2_0_targ_ht_axi_m_arburst),
        .o_l2_0_targ_ht_axi_m_arcache(o_l2_0_targ_ht_axi_m_arcache),
        .o_l2_0_targ_ht_axi_m_arid(o_l2_0_targ_ht_axi_m_arid),
        .o_l2_0_targ_ht_axi_m_arlen(o_l2_0_targ_ht_axi_m_arlen),
        .o_l2_0_targ_ht_axi_m_arlock(o_l2_0_targ_ht_axi_m_arlock),
        .o_l2_0_targ_ht_axi_m_arprot(o_l2_0_targ_ht_axi_m_arprot),
        .i_l2_0_targ_ht_axi_m_arready(i_l2_0_targ_ht_axi_m_arready),
        .o_l2_0_targ_ht_axi_m_arsize(o_l2_0_targ_ht_axi_m_arsize),
        .o_l2_0_targ_ht_axi_m_arvalid(o_l2_0_targ_ht_axi_m_arvalid),
        .i_l2_0_targ_ht_axi_m_rdata(i_l2_0_targ_ht_axi_m_rdata),
        .i_l2_0_targ_ht_axi_m_rid(i_l2_0_targ_ht_axi_m_rid),
        .i_l2_0_targ_ht_axi_m_rlast(i_l2_0_targ_ht_axi_m_rlast),
        .o_l2_0_targ_ht_axi_m_rready(o_l2_0_targ_ht_axi_m_rready),
        .i_l2_0_targ_ht_axi_m_rresp(i_l2_0_targ_ht_axi_m_rresp),
        .i_l2_0_targ_ht_axi_m_rvalid(i_l2_0_targ_ht_axi_m_rvalid),
        .o_l2_0_targ_ht_axi_m_awaddr(o_l2_0_targ_ht_axi_m_awaddr),
        .o_l2_0_targ_ht_axi_m_awburst(o_l2_0_targ_ht_axi_m_awburst),
        .o_l2_0_targ_ht_axi_m_awcache(o_l2_0_targ_ht_axi_m_awcache),
        .o_l2_0_targ_ht_axi_m_awid(o_l2_0_targ_ht_axi_m_awid),
        .o_l2_0_targ_ht_axi_m_awlen(o_l2_0_targ_ht_axi_m_awlen),
        .o_l2_0_targ_ht_axi_m_awlock(o_l2_0_targ_ht_axi_m_awlock),
        .o_l2_0_targ_ht_axi_m_awprot(o_l2_0_targ_ht_axi_m_awprot),
        .i_l2_0_targ_ht_axi_m_awready(i_l2_0_targ_ht_axi_m_awready),
        .o_l2_0_targ_ht_axi_m_awsize(o_l2_0_targ_ht_axi_m_awsize),
        .o_l2_0_targ_ht_axi_m_awvalid(o_l2_0_targ_ht_axi_m_awvalid),
        .i_l2_0_targ_ht_axi_m_bid(i_l2_0_targ_ht_axi_m_bid),
        .o_l2_0_targ_ht_axi_m_bready(o_l2_0_targ_ht_axi_m_bready),
        .i_l2_0_targ_ht_axi_m_bresp(i_l2_0_targ_ht_axi_m_bresp),
        .i_l2_0_targ_ht_axi_m_bvalid(i_l2_0_targ_ht_axi_m_bvalid),
        .o_l2_0_targ_ht_axi_m_wdata(o_l2_0_targ_ht_axi_m_wdata),
        .o_l2_0_targ_ht_axi_m_wlast(o_l2_0_targ_ht_axi_m_wlast),
        .i_l2_0_targ_ht_axi_m_wready(i_l2_0_targ_ht_axi_m_wready),
        .o_l2_0_targ_ht_axi_m_wstrb(o_l2_0_targ_ht_axi_m_wstrb),
        .o_l2_0_targ_ht_axi_m_wvalid(o_l2_0_targ_ht_axi_m_wvalid),
        .o_l2_0_targ_syscfg_apb_m_paddr(o_l2_0_targ_syscfg_apb_m_paddr),
        .o_l2_0_targ_syscfg_apb_m_penable(o_l2_0_targ_syscfg_apb_m_penable),
        .o_l2_0_targ_syscfg_apb_m_pprot(o_l2_0_targ_syscfg_apb_m_pprot),
        .i_l2_0_targ_syscfg_apb_m_prdata(i_l2_0_targ_syscfg_apb_m_prdata),
        .i_l2_0_targ_syscfg_apb_m_pready(i_l2_0_targ_syscfg_apb_m_pready),
        .o_l2_0_targ_syscfg_apb_m_psel(o_l2_0_targ_syscfg_apb_m_psel),
        .i_l2_0_targ_syscfg_apb_m_pslverr(i_l2_0_targ_syscfg_apb_m_pslverr),
        .o_l2_0_targ_syscfg_apb_m_pstrb(o_l2_0_targ_syscfg_apb_m_pstrb),
        .o_l2_0_targ_syscfg_apb_m_pwdata(o_l2_0_targ_syscfg_apb_m_pwdata),
        .o_l2_0_targ_syscfg_apb_m_pwrite(o_l2_0_targ_syscfg_apb_m_pwrite),
        .i_l2_1_aon_clk(i_l2_1_aon_clk),
        .i_l2_1_aon_rst_n(i_l2_1_aon_rst_n),
        .i_l2_1_clk(i_l2_1_clk),
        .i_l2_1_clken(i_l2_1_clken),
        .o_l2_1_pwr_idle_val(o_l2_1_pwr_idle_val),
        .o_l2_1_pwr_idle_ack(o_l2_1_pwr_idle_ack),
        .i_l2_1_pwr_idle_req(i_l2_1_pwr_idle_req),
        .i_l2_1_rst_n(i_l2_1_rst_n),
        .o_l2_1_targ_ht_axi_m_araddr(o_l2_1_targ_ht_axi_m_araddr),
        .o_l2_1_targ_ht_axi_m_arburst(o_l2_1_targ_ht_axi_m_arburst),
        .o_l2_1_targ_ht_axi_m_arcache(o_l2_1_targ_ht_axi_m_arcache),
        .o_l2_1_targ_ht_axi_m_arid(o_l2_1_targ_ht_axi_m_arid),
        .o_l2_1_targ_ht_axi_m_arlen(o_l2_1_targ_ht_axi_m_arlen),
        .o_l2_1_targ_ht_axi_m_arlock(o_l2_1_targ_ht_axi_m_arlock),
        .o_l2_1_targ_ht_axi_m_arprot(o_l2_1_targ_ht_axi_m_arprot),
        .i_l2_1_targ_ht_axi_m_arready(i_l2_1_targ_ht_axi_m_arready),
        .o_l2_1_targ_ht_axi_m_arsize(o_l2_1_targ_ht_axi_m_arsize),
        .o_l2_1_targ_ht_axi_m_arvalid(o_l2_1_targ_ht_axi_m_arvalid),
        .i_l2_1_targ_ht_axi_m_rdata(i_l2_1_targ_ht_axi_m_rdata),
        .i_l2_1_targ_ht_axi_m_rid(i_l2_1_targ_ht_axi_m_rid),
        .i_l2_1_targ_ht_axi_m_rlast(i_l2_1_targ_ht_axi_m_rlast),
        .o_l2_1_targ_ht_axi_m_rready(o_l2_1_targ_ht_axi_m_rready),
        .i_l2_1_targ_ht_axi_m_rresp(i_l2_1_targ_ht_axi_m_rresp),
        .i_l2_1_targ_ht_axi_m_rvalid(i_l2_1_targ_ht_axi_m_rvalid),
        .o_l2_1_targ_ht_axi_m_awaddr(o_l2_1_targ_ht_axi_m_awaddr),
        .o_l2_1_targ_ht_axi_m_awburst(o_l2_1_targ_ht_axi_m_awburst),
        .o_l2_1_targ_ht_axi_m_awcache(o_l2_1_targ_ht_axi_m_awcache),
        .o_l2_1_targ_ht_axi_m_awid(o_l2_1_targ_ht_axi_m_awid),
        .o_l2_1_targ_ht_axi_m_awlen(o_l2_1_targ_ht_axi_m_awlen),
        .o_l2_1_targ_ht_axi_m_awlock(o_l2_1_targ_ht_axi_m_awlock),
        .o_l2_1_targ_ht_axi_m_awprot(o_l2_1_targ_ht_axi_m_awprot),
        .i_l2_1_targ_ht_axi_m_awready(i_l2_1_targ_ht_axi_m_awready),
        .o_l2_1_targ_ht_axi_m_awsize(o_l2_1_targ_ht_axi_m_awsize),
        .o_l2_1_targ_ht_axi_m_awvalid(o_l2_1_targ_ht_axi_m_awvalid),
        .i_l2_1_targ_ht_axi_m_bid(i_l2_1_targ_ht_axi_m_bid),
        .o_l2_1_targ_ht_axi_m_bready(o_l2_1_targ_ht_axi_m_bready),
        .i_l2_1_targ_ht_axi_m_bresp(i_l2_1_targ_ht_axi_m_bresp),
        .i_l2_1_targ_ht_axi_m_bvalid(i_l2_1_targ_ht_axi_m_bvalid),
        .o_l2_1_targ_ht_axi_m_wdata(o_l2_1_targ_ht_axi_m_wdata),
        .o_l2_1_targ_ht_axi_m_wlast(o_l2_1_targ_ht_axi_m_wlast),
        .i_l2_1_targ_ht_axi_m_wready(i_l2_1_targ_ht_axi_m_wready),
        .o_l2_1_targ_ht_axi_m_wstrb(o_l2_1_targ_ht_axi_m_wstrb),
        .o_l2_1_targ_ht_axi_m_wvalid(o_l2_1_targ_ht_axi_m_wvalid),
        .o_l2_1_targ_syscfg_apb_m_paddr(o_l2_1_targ_syscfg_apb_m_paddr),
        .o_l2_1_targ_syscfg_apb_m_penable(o_l2_1_targ_syscfg_apb_m_penable),
        .o_l2_1_targ_syscfg_apb_m_pprot(o_l2_1_targ_syscfg_apb_m_pprot),
        .i_l2_1_targ_syscfg_apb_m_prdata(i_l2_1_targ_syscfg_apb_m_prdata),
        .i_l2_1_targ_syscfg_apb_m_pready(i_l2_1_targ_syscfg_apb_m_pready),
        .o_l2_1_targ_syscfg_apb_m_psel(o_l2_1_targ_syscfg_apb_m_psel),
        .i_l2_1_targ_syscfg_apb_m_pslverr(i_l2_1_targ_syscfg_apb_m_pslverr),
        .o_l2_1_targ_syscfg_apb_m_pstrb(o_l2_1_targ_syscfg_apb_m_pstrb),
        .o_l2_1_targ_syscfg_apb_m_pwdata(o_l2_1_targ_syscfg_apb_m_pwdata),
        .o_l2_1_targ_syscfg_apb_m_pwrite(o_l2_1_targ_syscfg_apb_m_pwrite),
        .i_l2_2_aon_clk(i_l2_2_aon_clk),
        .i_l2_2_aon_rst_n(i_l2_2_aon_rst_n),
        .i_l2_2_clk(i_l2_2_clk),
        .i_l2_2_clken(i_l2_2_clken),
        .o_l2_2_pwr_idle_val(o_l2_2_pwr_idle_val),
        .o_l2_2_pwr_idle_ack(o_l2_2_pwr_idle_ack),
        .i_l2_2_pwr_idle_req(i_l2_2_pwr_idle_req),
        .i_l2_2_rst_n(i_l2_2_rst_n),
        .o_l2_2_targ_ht_axi_m_araddr(o_l2_2_targ_ht_axi_m_araddr),
        .o_l2_2_targ_ht_axi_m_arburst(o_l2_2_targ_ht_axi_m_arburst),
        .o_l2_2_targ_ht_axi_m_arcache(o_l2_2_targ_ht_axi_m_arcache),
        .o_l2_2_targ_ht_axi_m_arid(o_l2_2_targ_ht_axi_m_arid),
        .o_l2_2_targ_ht_axi_m_arlen(o_l2_2_targ_ht_axi_m_arlen),
        .o_l2_2_targ_ht_axi_m_arlock(o_l2_2_targ_ht_axi_m_arlock),
        .o_l2_2_targ_ht_axi_m_arprot(o_l2_2_targ_ht_axi_m_arprot),
        .i_l2_2_targ_ht_axi_m_arready(i_l2_2_targ_ht_axi_m_arready),
        .o_l2_2_targ_ht_axi_m_arsize(o_l2_2_targ_ht_axi_m_arsize),
        .o_l2_2_targ_ht_axi_m_arvalid(o_l2_2_targ_ht_axi_m_arvalid),
        .i_l2_2_targ_ht_axi_m_rdata(i_l2_2_targ_ht_axi_m_rdata),
        .i_l2_2_targ_ht_axi_m_rid(i_l2_2_targ_ht_axi_m_rid),
        .i_l2_2_targ_ht_axi_m_rlast(i_l2_2_targ_ht_axi_m_rlast),
        .o_l2_2_targ_ht_axi_m_rready(o_l2_2_targ_ht_axi_m_rready),
        .i_l2_2_targ_ht_axi_m_rresp(i_l2_2_targ_ht_axi_m_rresp),
        .i_l2_2_targ_ht_axi_m_rvalid(i_l2_2_targ_ht_axi_m_rvalid),
        .o_l2_2_targ_ht_axi_m_awaddr(o_l2_2_targ_ht_axi_m_awaddr),
        .o_l2_2_targ_ht_axi_m_awburst(o_l2_2_targ_ht_axi_m_awburst),
        .o_l2_2_targ_ht_axi_m_awcache(o_l2_2_targ_ht_axi_m_awcache),
        .o_l2_2_targ_ht_axi_m_awid(o_l2_2_targ_ht_axi_m_awid),
        .o_l2_2_targ_ht_axi_m_awlen(o_l2_2_targ_ht_axi_m_awlen),
        .o_l2_2_targ_ht_axi_m_awlock(o_l2_2_targ_ht_axi_m_awlock),
        .o_l2_2_targ_ht_axi_m_awprot(o_l2_2_targ_ht_axi_m_awprot),
        .i_l2_2_targ_ht_axi_m_awready(i_l2_2_targ_ht_axi_m_awready),
        .o_l2_2_targ_ht_axi_m_awsize(o_l2_2_targ_ht_axi_m_awsize),
        .o_l2_2_targ_ht_axi_m_awvalid(o_l2_2_targ_ht_axi_m_awvalid),
        .i_l2_2_targ_ht_axi_m_bid(i_l2_2_targ_ht_axi_m_bid),
        .o_l2_2_targ_ht_axi_m_bready(o_l2_2_targ_ht_axi_m_bready),
        .i_l2_2_targ_ht_axi_m_bresp(i_l2_2_targ_ht_axi_m_bresp),
        .i_l2_2_targ_ht_axi_m_bvalid(i_l2_2_targ_ht_axi_m_bvalid),
        .o_l2_2_targ_ht_axi_m_wdata(o_l2_2_targ_ht_axi_m_wdata),
        .o_l2_2_targ_ht_axi_m_wlast(o_l2_2_targ_ht_axi_m_wlast),
        .i_l2_2_targ_ht_axi_m_wready(i_l2_2_targ_ht_axi_m_wready),
        .o_l2_2_targ_ht_axi_m_wstrb(o_l2_2_targ_ht_axi_m_wstrb),
        .o_l2_2_targ_ht_axi_m_wvalid(o_l2_2_targ_ht_axi_m_wvalid),
        .o_l2_2_targ_syscfg_apb_m_paddr(o_l2_2_targ_syscfg_apb_m_paddr),
        .o_l2_2_targ_syscfg_apb_m_penable(o_l2_2_targ_syscfg_apb_m_penable),
        .o_l2_2_targ_syscfg_apb_m_pprot(o_l2_2_targ_syscfg_apb_m_pprot),
        .i_l2_2_targ_syscfg_apb_m_prdata(i_l2_2_targ_syscfg_apb_m_prdata),
        .i_l2_2_targ_syscfg_apb_m_pready(i_l2_2_targ_syscfg_apb_m_pready),
        .o_l2_2_targ_syscfg_apb_m_psel(o_l2_2_targ_syscfg_apb_m_psel),
        .i_l2_2_targ_syscfg_apb_m_pslverr(i_l2_2_targ_syscfg_apb_m_pslverr),
        .o_l2_2_targ_syscfg_apb_m_pstrb(o_l2_2_targ_syscfg_apb_m_pstrb),
        .o_l2_2_targ_syscfg_apb_m_pwdata(o_l2_2_targ_syscfg_apb_m_pwdata),
        .o_l2_2_targ_syscfg_apb_m_pwrite(o_l2_2_targ_syscfg_apb_m_pwrite),
        .i_l2_3_aon_clk(i_l2_3_aon_clk),
        .i_l2_3_aon_rst_n(i_l2_3_aon_rst_n),
        .i_l2_3_clk(i_l2_3_clk),
        .i_l2_3_clken(i_l2_3_clken),
        .o_l2_3_pwr_idle_val(o_l2_3_pwr_idle_val),
        .o_l2_3_pwr_idle_ack(o_l2_3_pwr_idle_ack),
        .i_l2_3_pwr_idle_req(i_l2_3_pwr_idle_req),
        .i_l2_3_rst_n(i_l2_3_rst_n),
        .o_l2_3_targ_ht_axi_m_araddr(o_l2_3_targ_ht_axi_m_araddr),
        .o_l2_3_targ_ht_axi_m_arburst(o_l2_3_targ_ht_axi_m_arburst),
        .o_l2_3_targ_ht_axi_m_arcache(o_l2_3_targ_ht_axi_m_arcache),
        .o_l2_3_targ_ht_axi_m_arid(o_l2_3_targ_ht_axi_m_arid),
        .o_l2_3_targ_ht_axi_m_arlen(o_l2_3_targ_ht_axi_m_arlen),
        .o_l2_3_targ_ht_axi_m_arlock(o_l2_3_targ_ht_axi_m_arlock),
        .o_l2_3_targ_ht_axi_m_arprot(o_l2_3_targ_ht_axi_m_arprot),
        .i_l2_3_targ_ht_axi_m_arready(i_l2_3_targ_ht_axi_m_arready),
        .o_l2_3_targ_ht_axi_m_arsize(o_l2_3_targ_ht_axi_m_arsize),
        .o_l2_3_targ_ht_axi_m_arvalid(o_l2_3_targ_ht_axi_m_arvalid),
        .i_l2_3_targ_ht_axi_m_rdata(i_l2_3_targ_ht_axi_m_rdata),
        .i_l2_3_targ_ht_axi_m_rid(i_l2_3_targ_ht_axi_m_rid),
        .i_l2_3_targ_ht_axi_m_rlast(i_l2_3_targ_ht_axi_m_rlast),
        .o_l2_3_targ_ht_axi_m_rready(o_l2_3_targ_ht_axi_m_rready),
        .i_l2_3_targ_ht_axi_m_rresp(i_l2_3_targ_ht_axi_m_rresp),
        .i_l2_3_targ_ht_axi_m_rvalid(i_l2_3_targ_ht_axi_m_rvalid),
        .o_l2_3_targ_ht_axi_m_awaddr(o_l2_3_targ_ht_axi_m_awaddr),
        .o_l2_3_targ_ht_axi_m_awburst(o_l2_3_targ_ht_axi_m_awburst),
        .o_l2_3_targ_ht_axi_m_awcache(o_l2_3_targ_ht_axi_m_awcache),
        .o_l2_3_targ_ht_axi_m_awid(o_l2_3_targ_ht_axi_m_awid),
        .o_l2_3_targ_ht_axi_m_awlen(o_l2_3_targ_ht_axi_m_awlen),
        .o_l2_3_targ_ht_axi_m_awlock(o_l2_3_targ_ht_axi_m_awlock),
        .o_l2_3_targ_ht_axi_m_awprot(o_l2_3_targ_ht_axi_m_awprot),
        .i_l2_3_targ_ht_axi_m_awready(i_l2_3_targ_ht_axi_m_awready),
        .o_l2_3_targ_ht_axi_m_awsize(o_l2_3_targ_ht_axi_m_awsize),
        .o_l2_3_targ_ht_axi_m_awvalid(o_l2_3_targ_ht_axi_m_awvalid),
        .i_l2_3_targ_ht_axi_m_bid(i_l2_3_targ_ht_axi_m_bid),
        .o_l2_3_targ_ht_axi_m_bready(o_l2_3_targ_ht_axi_m_bready),
        .i_l2_3_targ_ht_axi_m_bresp(i_l2_3_targ_ht_axi_m_bresp),
        .i_l2_3_targ_ht_axi_m_bvalid(i_l2_3_targ_ht_axi_m_bvalid),
        .o_l2_3_targ_ht_axi_m_wdata(o_l2_3_targ_ht_axi_m_wdata),
        .o_l2_3_targ_ht_axi_m_wlast(o_l2_3_targ_ht_axi_m_wlast),
        .i_l2_3_targ_ht_axi_m_wready(i_l2_3_targ_ht_axi_m_wready),
        .o_l2_3_targ_ht_axi_m_wstrb(o_l2_3_targ_ht_axi_m_wstrb),
        .o_l2_3_targ_ht_axi_m_wvalid(o_l2_3_targ_ht_axi_m_wvalid),
        .o_l2_3_targ_syscfg_apb_m_paddr(o_l2_3_targ_syscfg_apb_m_paddr),
        .o_l2_3_targ_syscfg_apb_m_penable(o_l2_3_targ_syscfg_apb_m_penable),
        .o_l2_3_targ_syscfg_apb_m_pprot(o_l2_3_targ_syscfg_apb_m_pprot),
        .i_l2_3_targ_syscfg_apb_m_prdata(i_l2_3_targ_syscfg_apb_m_prdata),
        .i_l2_3_targ_syscfg_apb_m_pready(i_l2_3_targ_syscfg_apb_m_pready),
        .o_l2_3_targ_syscfg_apb_m_psel(o_l2_3_targ_syscfg_apb_m_psel),
        .i_l2_3_targ_syscfg_apb_m_pslverr(i_l2_3_targ_syscfg_apb_m_pslverr),
        .o_l2_3_targ_syscfg_apb_m_pstrb(o_l2_3_targ_syscfg_apb_m_pstrb),
        .o_l2_3_targ_syscfg_apb_m_pwdata(o_l2_3_targ_syscfg_apb_m_pwdata),
        .o_l2_3_targ_syscfg_apb_m_pwrite(o_l2_3_targ_syscfg_apb_m_pwrite),
        .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
        .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
        .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
        .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
        .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
        .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
        .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
        .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
        .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
        .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
        .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
        .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),

        // Token Network IOs
        // - Fences
        .o_aic_0_pwr_tok_idle_val(o_aic_0_pwr_tok_idle_val),
        .o_aic_0_pwr_tok_idle_ack(o_aic_0_pwr_tok_idle_ack),
        .i_aic_0_pwr_tok_idle_req(i_aic_0_pwr_tok_idle_req),
        .o_aic_1_pwr_tok_idle_val(o_aic_1_pwr_tok_idle_val),
        .o_aic_1_pwr_tok_idle_ack(o_aic_1_pwr_tok_idle_ack),
        .i_aic_1_pwr_tok_idle_req(i_aic_1_pwr_tok_idle_req),
        .o_aic_2_pwr_tok_idle_val(o_aic_2_pwr_tok_idle_val),
        .o_aic_2_pwr_tok_idle_ack(o_aic_2_pwr_tok_idle_ack),
        .i_aic_2_pwr_tok_idle_req(i_aic_2_pwr_tok_idle_req),
        .o_aic_3_pwr_tok_idle_val(o_aic_3_pwr_tok_idle_val),
        .o_aic_3_pwr_tok_idle_ack(o_aic_3_pwr_tok_idle_ack),
        .i_aic_3_pwr_tok_idle_req(i_aic_3_pwr_tok_idle_req),

        // - NIUs
        .i_aic_0_init_tok_ocpl_s_maddr(i_aic_0_init_tok_ocpl_s_maddr),
        .i_aic_0_init_tok_ocpl_s_mcmd(i_aic_0_init_tok_ocpl_s_mcmd),
        .i_aic_0_init_tok_ocpl_s_mdata(i_aic_0_init_tok_ocpl_s_mdata),
        .o_aic_0_init_tok_ocpl_s_scmdaccept(o_aic_0_init_tok_ocpl_s_scmdaccept),
        .o_aic_0_targ_tok_ocpl_m_maddr(o_aic_0_targ_tok_ocpl_m_maddr),
        .o_aic_0_targ_tok_ocpl_m_mcmd(o_aic_0_targ_tok_ocpl_m_mcmd),
        .o_aic_0_targ_tok_ocpl_m_mdata(o_aic_0_targ_tok_ocpl_m_mdata),
        .i_aic_0_targ_tok_ocpl_m_scmdaccept(i_aic_0_targ_tok_ocpl_m_scmdaccept),
        .i_aic_1_init_tok_ocpl_s_maddr(i_aic_1_init_tok_ocpl_s_maddr),
        .i_aic_1_init_tok_ocpl_s_mcmd(i_aic_1_init_tok_ocpl_s_mcmd),
        .i_aic_1_init_tok_ocpl_s_mdata(i_aic_1_init_tok_ocpl_s_mdata),
        .o_aic_1_init_tok_ocpl_s_scmdaccept(o_aic_1_init_tok_ocpl_s_scmdaccept),
        .o_aic_1_targ_tok_ocpl_m_maddr(o_aic_1_targ_tok_ocpl_m_maddr),
        .o_aic_1_targ_tok_ocpl_m_mcmd(o_aic_1_targ_tok_ocpl_m_mcmd),
        .o_aic_1_targ_tok_ocpl_m_mdata(o_aic_1_targ_tok_ocpl_m_mdata),
        .i_aic_1_targ_tok_ocpl_m_scmdaccept(i_aic_1_targ_tok_ocpl_m_scmdaccept),
        .i_aic_2_init_tok_ocpl_s_maddr(i_aic_2_init_tok_ocpl_s_maddr),
        .i_aic_2_init_tok_ocpl_s_mcmd(i_aic_2_init_tok_ocpl_s_mcmd),
        .i_aic_2_init_tok_ocpl_s_mdata(i_aic_2_init_tok_ocpl_s_mdata),
        .o_aic_2_init_tok_ocpl_s_scmdaccept(o_aic_2_init_tok_ocpl_s_scmdaccept),
        .o_aic_2_targ_tok_ocpl_m_maddr(o_aic_2_targ_tok_ocpl_m_maddr),
        .o_aic_2_targ_tok_ocpl_m_mcmd(o_aic_2_targ_tok_ocpl_m_mcmd),
        .o_aic_2_targ_tok_ocpl_m_mdata(o_aic_2_targ_tok_ocpl_m_mdata),
        .i_aic_2_targ_tok_ocpl_m_scmdaccept(i_aic_2_targ_tok_ocpl_m_scmdaccept),
        .o_aic_3_targ_tok_ocpl_m_maddr(o_aic_3_targ_tok_ocpl_m_maddr),
        .o_aic_3_targ_tok_ocpl_m_mcmd(o_aic_3_targ_tok_ocpl_m_mcmd),
        .o_aic_3_targ_tok_ocpl_m_mdata(o_aic_3_targ_tok_ocpl_m_mdata),
        .i_aic_3_targ_tok_ocpl_m_scmdaccept(i_aic_3_targ_tok_ocpl_m_scmdaccept),
        .i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data),
        .i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head),
        .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy),
        .i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail),
        .i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld),
        .i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data),
        .i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head),
        .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy),
        .i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail),
        .i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld),
        .o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data),
        .o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head),
        .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy),
        .o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail),
        .o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld),
        .o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data),
        .o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head),
        .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy),
        .o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail),
        .o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld),

        .i_noc_clk(i_noc_clk),
        .i_noc_rst_n(i_noc_rst_n),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  )
    );

    // Instance of noc_h_west_p
    noc_h_west_p h_west_p (
        .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data),
        .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head),
        .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy),
        .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail),
        .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld),
        .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data),
        .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head),
        .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy),
        .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail),
        .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld),
        .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data),
        .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head),
        .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy),
        .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail),
        .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld),
        .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data),
        .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head),
        .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy),
        .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail),
        .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld),
        .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data),
        .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head),
        .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy),
        .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail),
        .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld),
        .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data),
        .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head),
        .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy),
        .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail),
        .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld),
        .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data),
        .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head),
        .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy),
        .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail),
        .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld),
        .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data),
        .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head),
        .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy),
        .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail),
        .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld),
        .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data),
        .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head),
        .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy),
        .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail),
        .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld),
        .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data),
        .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head),
        .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy),
        .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail),
        .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld),
        .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_data),
        .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_head),
        .i_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_rdy),
        .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_tail),
        .o_dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld(dp_lnk_cross_west_to_ddrw_256_0_egr_to_lnk_cross_west_to_ddrw_256_0_ingr_vld),
        .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_data),
        .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_head),
        .o_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_rdy),
        .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_tail),
        .i_dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld(dp_lnk_cross_west_to_ddrw_256_0_ingr_resp_to_lnk_cross_west_to_ddrw_256_0_egr_resp_vld),
        .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_data),
        .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_head),
        .i_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_rdy),
        .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_tail),
        .o_dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld(dp_lnk_cross_west_to_ddrw_256_1_egr_to_lnk_cross_west_to_ddrw_256_1_ingr_vld),
        .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_data),
        .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_head),
        .o_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_rdy),
        .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_tail),
        .i_dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld(dp_lnk_cross_west_to_ddrw_256_1_ingr_resp_to_lnk_cross_west_to_ddrw_256_1_egr_resp_vld),
        .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_data),
        .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_head),
        .i_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_rdy),
        .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_tail),
        .o_dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld(dp_lnk_cross_west_to_ddrw_256_2_egr_to_lnk_cross_west_to_ddrw_256_2_ingr_vld),
        .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_data),
        .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_head),
        .o_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_rdy),
        .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_tail),
        .i_dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld(dp_lnk_cross_west_to_ddrw_256_2_ingr_resp_to_lnk_cross_west_to_ddrw_256_2_egr_resp_vld),
        .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_data),
        .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_head),
        .i_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_rdy),
        .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_tail),
        .o_dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld(dp_lnk_cross_west_to_ddrw_256_3_egr_to_lnk_cross_west_to_ddrw_256_3_ingr_vld),
        .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_data),
        .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_head),
        .o_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_rdy),
        .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_tail),
        .i_dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld(dp_lnk_cross_west_to_ddrw_256_3_ingr_resp_to_lnk_cross_west_to_ddrw_256_3_egr_resp_vld),
        .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_data),
        .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_head),
        .i_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_rdy),
        .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_tail),
        .o_dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld(dp_lnk_cross_west_to_ddrw_32_egr_to_lnk_cross_west_to_ddrw_32_ingr_vld),
        .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_data),
        .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_head),
        .o_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_rdy),
        .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_tail),
        .i_dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld(dp_lnk_cross_west_to_ddrw_32_ingr_resp_to_lnk_cross_west_to_ddrw_32_egr_resp_vld),
        .i_noc_clk(i_noc_clk),
        .i_noc_rst_n(i_noc_rst_n),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  ),
        .bisr_clk('0),
        .bisr_reset('0),
        .bisr_shift_en('0),
        .bisr_si('0),
        .bisr_so(  )
    );

    // Instance of noc_soc_p
    noc_soc_p soc_p (
        .i_apu_aon_clk(i_apu_aon_clk),
        .i_apu_aon_rst_n(i_apu_aon_rst_n),
        .i_apu_init_lt_axi_s_araddr(i_apu_init_lt_axi_s_araddr),
        .i_apu_init_lt_axi_s_arburst(i_apu_init_lt_axi_s_arburst),
        .i_apu_init_lt_axi_s_arcache(i_apu_init_lt_axi_s_arcache),
        .i_apu_init_lt_axi_s_arid(i_apu_init_lt_axi_s_arid),
        .i_apu_init_lt_axi_s_arlen(i_apu_init_lt_axi_s_arlen),
        .i_apu_init_lt_axi_s_arlock(i_apu_init_lt_axi_s_arlock),
        .i_apu_init_lt_axi_s_arprot(i_apu_init_lt_axi_s_arprot),
        .i_apu_init_lt_axi_s_arqos(i_apu_init_lt_axi_s_arqos),
        .o_apu_init_lt_axi_s_arready(o_apu_init_lt_axi_s_arready),
        .i_apu_init_lt_axi_s_arsize(i_apu_init_lt_axi_s_arsize),
        .i_apu_init_lt_axi_s_arvalid(i_apu_init_lt_axi_s_arvalid),
        .i_apu_init_lt_axi_s_awaddr(i_apu_init_lt_axi_s_awaddr),
        .i_apu_init_lt_axi_s_awburst(i_apu_init_lt_axi_s_awburst),
        .i_apu_init_lt_axi_s_awcache(i_apu_init_lt_axi_s_awcache),
        .i_apu_init_lt_axi_s_awid(i_apu_init_lt_axi_s_awid),
        .i_apu_init_lt_axi_s_awlen(i_apu_init_lt_axi_s_awlen),
        .i_apu_init_lt_axi_s_awlock(i_apu_init_lt_axi_s_awlock),
        .i_apu_init_lt_axi_s_awprot(i_apu_init_lt_axi_s_awprot),
        .i_apu_init_lt_axi_s_awqos(i_apu_init_lt_axi_s_awqos),
        .o_apu_init_lt_axi_s_awready(o_apu_init_lt_axi_s_awready),
        .i_apu_init_lt_axi_s_awsize(i_apu_init_lt_axi_s_awsize),
        .i_apu_init_lt_axi_s_awvalid(i_apu_init_lt_axi_s_awvalid),
        .o_apu_init_lt_axi_s_bid(o_apu_init_lt_axi_s_bid),
        .i_apu_init_lt_axi_s_bready(i_apu_init_lt_axi_s_bready),
        .o_apu_init_lt_axi_s_bresp(o_apu_init_lt_axi_s_bresp),
        .o_apu_init_lt_axi_s_bvalid(o_apu_init_lt_axi_s_bvalid),
        .o_apu_init_lt_axi_s_rdata(o_apu_init_lt_axi_s_rdata),
        .o_apu_init_lt_axi_s_rid(o_apu_init_lt_axi_s_rid),
        .o_apu_init_lt_axi_s_rlast(o_apu_init_lt_axi_s_rlast),
        .i_apu_init_lt_axi_s_rready(i_apu_init_lt_axi_s_rready),
        .o_apu_init_lt_axi_s_rresp(o_apu_init_lt_axi_s_rresp),
        .o_apu_init_lt_axi_s_rvalid(o_apu_init_lt_axi_s_rvalid),
        .i_apu_init_lt_axi_s_wdata(i_apu_init_lt_axi_s_wdata),
        .i_apu_init_lt_axi_s_wlast(i_apu_init_lt_axi_s_wlast),
        .o_apu_init_lt_axi_s_wready(o_apu_init_lt_axi_s_wready),
        .i_apu_init_lt_axi_s_wstrb(i_apu_init_lt_axi_s_wstrb),
        .i_apu_init_lt_axi_s_wvalid(i_apu_init_lt_axi_s_wvalid),
        .i_apu_init_mt_axi_s_araddr(i_apu_init_mt_axi_s_araddr),
        .i_apu_init_mt_axi_s_arburst(i_apu_init_mt_axi_s_arburst),
        .i_apu_init_mt_axi_s_arcache(i_apu_init_mt_axi_s_arcache),
        .i_apu_init_mt_axi_s_arid(i_apu_init_mt_axi_s_arid),
        .i_apu_init_mt_axi_s_arlen(i_apu_init_mt_axi_s_arlen),
        .i_apu_init_mt_axi_s_arlock(i_apu_init_mt_axi_s_arlock),
        .i_apu_init_mt_axi_s_arprot(i_apu_init_mt_axi_s_arprot),
        .i_apu_init_mt_axi_s_arqos(i_apu_init_mt_axi_s_arqos),
        .o_apu_init_mt_axi_s_arready(o_apu_init_mt_axi_s_arready),
        .i_apu_init_mt_axi_s_arsize(i_apu_init_mt_axi_s_arsize),
        .i_apu_init_mt_axi_s_arvalid(i_apu_init_mt_axi_s_arvalid),
        .o_apu_init_mt_axi_s_rdata(o_apu_init_mt_axi_s_rdata),
        .o_apu_init_mt_axi_s_rid(o_apu_init_mt_axi_s_rid),
        .o_apu_init_mt_axi_s_rlast(o_apu_init_mt_axi_s_rlast),
        .i_apu_init_mt_axi_s_rready(i_apu_init_mt_axi_s_rready),
        .o_apu_init_mt_axi_s_rresp(o_apu_init_mt_axi_s_rresp),
        .o_apu_init_mt_axi_s_rvalid(o_apu_init_mt_axi_s_rvalid),
        .i_apu_init_mt_axi_s_awaddr(i_apu_init_mt_axi_s_awaddr),
        .i_apu_init_mt_axi_s_awburst(i_apu_init_mt_axi_s_awburst),
        .i_apu_init_mt_axi_s_awcache(i_apu_init_mt_axi_s_awcache),
        .i_apu_init_mt_axi_s_awid(i_apu_init_mt_axi_s_awid),
        .i_apu_init_mt_axi_s_awlen(i_apu_init_mt_axi_s_awlen),
        .i_apu_init_mt_axi_s_awlock(i_apu_init_mt_axi_s_awlock),
        .i_apu_init_mt_axi_s_awprot(i_apu_init_mt_axi_s_awprot),
        .i_apu_init_mt_axi_s_awqos(i_apu_init_mt_axi_s_awqos),
        .o_apu_init_mt_axi_s_awready(o_apu_init_mt_axi_s_awready),
        .i_apu_init_mt_axi_s_awsize(i_apu_init_mt_axi_s_awsize),
        .i_apu_init_mt_axi_s_awvalid(i_apu_init_mt_axi_s_awvalid),
        .o_apu_init_mt_axi_s_bid(o_apu_init_mt_axi_s_bid),
        .i_apu_init_mt_axi_s_bready(i_apu_init_mt_axi_s_bready),
        .o_apu_init_mt_axi_s_bresp(o_apu_init_mt_axi_s_bresp),
        .o_apu_init_mt_axi_s_bvalid(o_apu_init_mt_axi_s_bvalid),
        .i_apu_init_mt_axi_s_wdata(i_apu_init_mt_axi_s_wdata),
        .i_apu_init_mt_axi_s_wlast(i_apu_init_mt_axi_s_wlast),
        .o_apu_init_mt_axi_s_wready(o_apu_init_mt_axi_s_wready),
        .i_apu_init_mt_axi_s_wstrb(i_apu_init_mt_axi_s_wstrb),
        .i_apu_init_mt_axi_s_wvalid(i_apu_init_mt_axi_s_wvalid),
        .o_apu_pwr_idle_val(o_apu_pwr_idle_val),
        .o_apu_pwr_idle_ack(o_apu_pwr_idle_ack),
        .i_apu_pwr_idle_req(i_apu_pwr_idle_req),
        .o_apu_targ_lt_axi_m_araddr(o_apu_targ_lt_axi_m_araddr),
        .o_apu_targ_lt_axi_m_arburst(o_apu_targ_lt_axi_m_arburst),
        .o_apu_targ_lt_axi_m_arcache(o_apu_targ_lt_axi_m_arcache),
        .o_apu_targ_lt_axi_m_arid(o_apu_targ_lt_axi_m_arid),
        .o_apu_targ_lt_axi_m_arlen(o_apu_targ_lt_axi_m_arlen),
        .o_apu_targ_lt_axi_m_arlock(o_apu_targ_lt_axi_m_arlock),
        .o_apu_targ_lt_axi_m_arprot(o_apu_targ_lt_axi_m_arprot),
        .o_apu_targ_lt_axi_m_arqos(o_apu_targ_lt_axi_m_arqos),
        .i_apu_targ_lt_axi_m_arready(i_apu_targ_lt_axi_m_arready),
        .o_apu_targ_lt_axi_m_arsize(o_apu_targ_lt_axi_m_arsize),
        .o_apu_targ_lt_axi_m_arvalid(o_apu_targ_lt_axi_m_arvalid),
        .o_apu_targ_lt_axi_m_awaddr(o_apu_targ_lt_axi_m_awaddr),
        .o_apu_targ_lt_axi_m_awburst(o_apu_targ_lt_axi_m_awburst),
        .o_apu_targ_lt_axi_m_awcache(o_apu_targ_lt_axi_m_awcache),
        .o_apu_targ_lt_axi_m_awid(o_apu_targ_lt_axi_m_awid),
        .o_apu_targ_lt_axi_m_awlen(o_apu_targ_lt_axi_m_awlen),
        .o_apu_targ_lt_axi_m_awlock(o_apu_targ_lt_axi_m_awlock),
        .o_apu_targ_lt_axi_m_awprot(o_apu_targ_lt_axi_m_awprot),
        .o_apu_targ_lt_axi_m_awqos(o_apu_targ_lt_axi_m_awqos),
        .i_apu_targ_lt_axi_m_awready(i_apu_targ_lt_axi_m_awready),
        .o_apu_targ_lt_axi_m_awsize(o_apu_targ_lt_axi_m_awsize),
        .o_apu_targ_lt_axi_m_awvalid(o_apu_targ_lt_axi_m_awvalid),
        .i_apu_targ_lt_axi_m_bid(i_apu_targ_lt_axi_m_bid),
        .o_apu_targ_lt_axi_m_bready(o_apu_targ_lt_axi_m_bready),
        .i_apu_targ_lt_axi_m_bresp(i_apu_targ_lt_axi_m_bresp),
        .i_apu_targ_lt_axi_m_bvalid(i_apu_targ_lt_axi_m_bvalid),
        .i_apu_targ_lt_axi_m_rdata(i_apu_targ_lt_axi_m_rdata),
        .i_apu_targ_lt_axi_m_rid(i_apu_targ_lt_axi_m_rid),
        .i_apu_targ_lt_axi_m_rlast(i_apu_targ_lt_axi_m_rlast),
        .o_apu_targ_lt_axi_m_rready(o_apu_targ_lt_axi_m_rready),
        .i_apu_targ_lt_axi_m_rresp(i_apu_targ_lt_axi_m_rresp),
        .i_apu_targ_lt_axi_m_rvalid(i_apu_targ_lt_axi_m_rvalid),
        .o_apu_targ_lt_axi_m_wdata(o_apu_targ_lt_axi_m_wdata),
        .o_apu_targ_lt_axi_m_wlast(o_apu_targ_lt_axi_m_wlast),
        .i_apu_targ_lt_axi_m_wready(i_apu_targ_lt_axi_m_wready),
        .o_apu_targ_lt_axi_m_wstrb(o_apu_targ_lt_axi_m_wstrb),
        .o_apu_targ_lt_axi_m_wvalid(o_apu_targ_lt_axi_m_wvalid),
        .o_apu_targ_syscfg_apb_m_paddr(o_apu_targ_syscfg_apb_m_paddr),
        .o_apu_targ_syscfg_apb_m_penable(o_apu_targ_syscfg_apb_m_penable),
        .o_apu_targ_syscfg_apb_m_pprot(o_apu_targ_syscfg_apb_m_pprot),
        .i_apu_targ_syscfg_apb_m_prdata(i_apu_targ_syscfg_apb_m_prdata),
        .i_apu_targ_syscfg_apb_m_pready(i_apu_targ_syscfg_apb_m_pready),
        .o_apu_targ_syscfg_apb_m_psel(o_apu_targ_syscfg_apb_m_psel),
        .i_apu_targ_syscfg_apb_m_pslverr(i_apu_targ_syscfg_apb_m_pslverr),
        .o_apu_targ_syscfg_apb_m_pstrb(o_apu_targ_syscfg_apb_m_pstrb),
        .o_apu_targ_syscfg_apb_m_pwdata(o_apu_targ_syscfg_apb_m_pwdata),
        .o_apu_targ_syscfg_apb_m_pwrite(o_apu_targ_syscfg_apb_m_pwrite),
        .i_apu_x_clk(i_apu_x_clk),
        .i_apu_x_clken(i_apu_x_clken),
        .i_apu_x_rst_n(i_apu_x_rst_n),
        .i_dcd_aon_clk(i_dcd_aon_clk),
        .i_dcd_aon_rst_n(i_dcd_aon_rst_n),
        .i_dcd_codec_clk(i_dcd_codec_clk),
        .i_dcd_codec_clken(i_dcd_codec_clken),
        .i_dcd_codec_rst_n(i_dcd_codec_rst_n),
        .i_dcd_dec_0_init_mt_axi_s_araddr(i_dcd_dec_0_init_mt_axi_s_araddr),
        .i_dcd_dec_0_init_mt_axi_s_arburst(i_dcd_dec_0_init_mt_axi_s_arburst),
        .i_dcd_dec_0_init_mt_axi_s_arcache(i_dcd_dec_0_init_mt_axi_s_arcache),
        .i_dcd_dec_0_init_mt_axi_s_arid(i_dcd_dec_0_init_mt_axi_s_arid),
        .i_dcd_dec_0_init_mt_axi_s_arlen(i_dcd_dec_0_init_mt_axi_s_arlen),
        .i_dcd_dec_0_init_mt_axi_s_arlock(i_dcd_dec_0_init_mt_axi_s_arlock),
        .i_dcd_dec_0_init_mt_axi_s_arprot(i_dcd_dec_0_init_mt_axi_s_arprot),
        .i_dcd_dec_0_init_mt_axi_s_arqos(i_dcd_dec_0_init_mt_axi_s_arqos),
        .o_dcd_dec_0_init_mt_axi_s_arready(o_dcd_dec_0_init_mt_axi_s_arready),
        .i_dcd_dec_0_init_mt_axi_s_arsize(i_dcd_dec_0_init_mt_axi_s_arsize),
        .i_dcd_dec_0_init_mt_axi_s_arvalid(i_dcd_dec_0_init_mt_axi_s_arvalid),
        .o_dcd_dec_0_init_mt_axi_s_rdata(o_dcd_dec_0_init_mt_axi_s_rdata),
        .o_dcd_dec_0_init_mt_axi_s_rid(o_dcd_dec_0_init_mt_axi_s_rid),
        .o_dcd_dec_0_init_mt_axi_s_rlast(o_dcd_dec_0_init_mt_axi_s_rlast),
        .i_dcd_dec_0_init_mt_axi_s_rready(i_dcd_dec_0_init_mt_axi_s_rready),
        .o_dcd_dec_0_init_mt_axi_s_rresp(o_dcd_dec_0_init_mt_axi_s_rresp),
        .o_dcd_dec_0_init_mt_axi_s_rvalid(o_dcd_dec_0_init_mt_axi_s_rvalid),
        .i_dcd_dec_0_init_mt_axi_s_awaddr(i_dcd_dec_0_init_mt_axi_s_awaddr),
        .i_dcd_dec_0_init_mt_axi_s_awburst(i_dcd_dec_0_init_mt_axi_s_awburst),
        .i_dcd_dec_0_init_mt_axi_s_awcache(i_dcd_dec_0_init_mt_axi_s_awcache),
        .i_dcd_dec_0_init_mt_axi_s_awid(i_dcd_dec_0_init_mt_axi_s_awid),
        .i_dcd_dec_0_init_mt_axi_s_awlen(i_dcd_dec_0_init_mt_axi_s_awlen),
        .i_dcd_dec_0_init_mt_axi_s_awlock(i_dcd_dec_0_init_mt_axi_s_awlock),
        .i_dcd_dec_0_init_mt_axi_s_awprot(i_dcd_dec_0_init_mt_axi_s_awprot),
        .i_dcd_dec_0_init_mt_axi_s_awqos(i_dcd_dec_0_init_mt_axi_s_awqos),
        .o_dcd_dec_0_init_mt_axi_s_awready(o_dcd_dec_0_init_mt_axi_s_awready),
        .i_dcd_dec_0_init_mt_axi_s_awsize(i_dcd_dec_0_init_mt_axi_s_awsize),
        .i_dcd_dec_0_init_mt_axi_s_awvalid(i_dcd_dec_0_init_mt_axi_s_awvalid),
        .o_dcd_dec_0_init_mt_axi_s_bid(o_dcd_dec_0_init_mt_axi_s_bid),
        .i_dcd_dec_0_init_mt_axi_s_bready(i_dcd_dec_0_init_mt_axi_s_bready),
        .o_dcd_dec_0_init_mt_axi_s_bresp(o_dcd_dec_0_init_mt_axi_s_bresp),
        .o_dcd_dec_0_init_mt_axi_s_bvalid(o_dcd_dec_0_init_mt_axi_s_bvalid),
        .i_dcd_dec_0_init_mt_axi_s_wdata(i_dcd_dec_0_init_mt_axi_s_wdata),
        .i_dcd_dec_0_init_mt_axi_s_wlast(i_dcd_dec_0_init_mt_axi_s_wlast),
        .o_dcd_dec_0_init_mt_axi_s_wready(o_dcd_dec_0_init_mt_axi_s_wready),
        .i_dcd_dec_0_init_mt_axi_s_wstrb(i_dcd_dec_0_init_mt_axi_s_wstrb),
        .i_dcd_dec_0_init_mt_axi_s_wvalid(i_dcd_dec_0_init_mt_axi_s_wvalid),
        .i_dcd_dec_1_init_mt_axi_s_araddr(i_dcd_dec_1_init_mt_axi_s_araddr),
        .i_dcd_dec_1_init_mt_axi_s_arburst(i_dcd_dec_1_init_mt_axi_s_arburst),
        .i_dcd_dec_1_init_mt_axi_s_arcache(i_dcd_dec_1_init_mt_axi_s_arcache),
        .i_dcd_dec_1_init_mt_axi_s_arid(i_dcd_dec_1_init_mt_axi_s_arid),
        .i_dcd_dec_1_init_mt_axi_s_arlen(i_dcd_dec_1_init_mt_axi_s_arlen),
        .i_dcd_dec_1_init_mt_axi_s_arlock(i_dcd_dec_1_init_mt_axi_s_arlock),
        .i_dcd_dec_1_init_mt_axi_s_arprot(i_dcd_dec_1_init_mt_axi_s_arprot),
        .i_dcd_dec_1_init_mt_axi_s_arqos(i_dcd_dec_1_init_mt_axi_s_arqos),
        .o_dcd_dec_1_init_mt_axi_s_arready(o_dcd_dec_1_init_mt_axi_s_arready),
        .i_dcd_dec_1_init_mt_axi_s_arsize(i_dcd_dec_1_init_mt_axi_s_arsize),
        .i_dcd_dec_1_init_mt_axi_s_arvalid(i_dcd_dec_1_init_mt_axi_s_arvalid),
        .o_dcd_dec_1_init_mt_axi_s_rdata(o_dcd_dec_1_init_mt_axi_s_rdata),
        .o_dcd_dec_1_init_mt_axi_s_rid(o_dcd_dec_1_init_mt_axi_s_rid),
        .o_dcd_dec_1_init_mt_axi_s_rlast(o_dcd_dec_1_init_mt_axi_s_rlast),
        .i_dcd_dec_1_init_mt_axi_s_rready(i_dcd_dec_1_init_mt_axi_s_rready),
        .o_dcd_dec_1_init_mt_axi_s_rresp(o_dcd_dec_1_init_mt_axi_s_rresp),
        .o_dcd_dec_1_init_mt_axi_s_rvalid(o_dcd_dec_1_init_mt_axi_s_rvalid),
        .i_dcd_dec_1_init_mt_axi_s_awaddr(i_dcd_dec_1_init_mt_axi_s_awaddr),
        .i_dcd_dec_1_init_mt_axi_s_awburst(i_dcd_dec_1_init_mt_axi_s_awburst),
        .i_dcd_dec_1_init_mt_axi_s_awcache(i_dcd_dec_1_init_mt_axi_s_awcache),
        .i_dcd_dec_1_init_mt_axi_s_awid(i_dcd_dec_1_init_mt_axi_s_awid),
        .i_dcd_dec_1_init_mt_axi_s_awlen(i_dcd_dec_1_init_mt_axi_s_awlen),
        .i_dcd_dec_1_init_mt_axi_s_awlock(i_dcd_dec_1_init_mt_axi_s_awlock),
        .i_dcd_dec_1_init_mt_axi_s_awprot(i_dcd_dec_1_init_mt_axi_s_awprot),
        .i_dcd_dec_1_init_mt_axi_s_awqos(i_dcd_dec_1_init_mt_axi_s_awqos),
        .o_dcd_dec_1_init_mt_axi_s_awready(o_dcd_dec_1_init_mt_axi_s_awready),
        .i_dcd_dec_1_init_mt_axi_s_awsize(i_dcd_dec_1_init_mt_axi_s_awsize),
        .i_dcd_dec_1_init_mt_axi_s_awvalid(i_dcd_dec_1_init_mt_axi_s_awvalid),
        .o_dcd_dec_1_init_mt_axi_s_bid(o_dcd_dec_1_init_mt_axi_s_bid),
        .i_dcd_dec_1_init_mt_axi_s_bready(i_dcd_dec_1_init_mt_axi_s_bready),
        .o_dcd_dec_1_init_mt_axi_s_bresp(o_dcd_dec_1_init_mt_axi_s_bresp),
        .o_dcd_dec_1_init_mt_axi_s_bvalid(o_dcd_dec_1_init_mt_axi_s_bvalid),
        .i_dcd_dec_1_init_mt_axi_s_wdata(i_dcd_dec_1_init_mt_axi_s_wdata),
        .i_dcd_dec_1_init_mt_axi_s_wlast(i_dcd_dec_1_init_mt_axi_s_wlast),
        .o_dcd_dec_1_init_mt_axi_s_wready(o_dcd_dec_1_init_mt_axi_s_wready),
        .i_dcd_dec_1_init_mt_axi_s_wstrb(i_dcd_dec_1_init_mt_axi_s_wstrb),
        .i_dcd_dec_1_init_mt_axi_s_wvalid(i_dcd_dec_1_init_mt_axi_s_wvalid),
        .i_dcd_dec_2_init_mt_axi_s_araddr(i_dcd_dec_2_init_mt_axi_s_araddr),
        .i_dcd_dec_2_init_mt_axi_s_arburst(i_dcd_dec_2_init_mt_axi_s_arburst),
        .i_dcd_dec_2_init_mt_axi_s_arcache(i_dcd_dec_2_init_mt_axi_s_arcache),
        .i_dcd_dec_2_init_mt_axi_s_arid(i_dcd_dec_2_init_mt_axi_s_arid),
        .i_dcd_dec_2_init_mt_axi_s_arlen(i_dcd_dec_2_init_mt_axi_s_arlen),
        .i_dcd_dec_2_init_mt_axi_s_arlock(i_dcd_dec_2_init_mt_axi_s_arlock),
        .i_dcd_dec_2_init_mt_axi_s_arprot(i_dcd_dec_2_init_mt_axi_s_arprot),
        .i_dcd_dec_2_init_mt_axi_s_arqos(i_dcd_dec_2_init_mt_axi_s_arqos),
        .o_dcd_dec_2_init_mt_axi_s_arready(o_dcd_dec_2_init_mt_axi_s_arready),
        .i_dcd_dec_2_init_mt_axi_s_arsize(i_dcd_dec_2_init_mt_axi_s_arsize),
        .i_dcd_dec_2_init_mt_axi_s_arvalid(i_dcd_dec_2_init_mt_axi_s_arvalid),
        .o_dcd_dec_2_init_mt_axi_s_rdata(o_dcd_dec_2_init_mt_axi_s_rdata),
        .o_dcd_dec_2_init_mt_axi_s_rid(o_dcd_dec_2_init_mt_axi_s_rid),
        .o_dcd_dec_2_init_mt_axi_s_rlast(o_dcd_dec_2_init_mt_axi_s_rlast),
        .i_dcd_dec_2_init_mt_axi_s_rready(i_dcd_dec_2_init_mt_axi_s_rready),
        .o_dcd_dec_2_init_mt_axi_s_rresp(o_dcd_dec_2_init_mt_axi_s_rresp),
        .o_dcd_dec_2_init_mt_axi_s_rvalid(o_dcd_dec_2_init_mt_axi_s_rvalid),
        .i_dcd_dec_2_init_mt_axi_s_awaddr(i_dcd_dec_2_init_mt_axi_s_awaddr),
        .i_dcd_dec_2_init_mt_axi_s_awburst(i_dcd_dec_2_init_mt_axi_s_awburst),
        .i_dcd_dec_2_init_mt_axi_s_awcache(i_dcd_dec_2_init_mt_axi_s_awcache),
        .i_dcd_dec_2_init_mt_axi_s_awid(i_dcd_dec_2_init_mt_axi_s_awid),
        .i_dcd_dec_2_init_mt_axi_s_awlen(i_dcd_dec_2_init_mt_axi_s_awlen),
        .i_dcd_dec_2_init_mt_axi_s_awlock(i_dcd_dec_2_init_mt_axi_s_awlock),
        .i_dcd_dec_2_init_mt_axi_s_awprot(i_dcd_dec_2_init_mt_axi_s_awprot),
        .i_dcd_dec_2_init_mt_axi_s_awqos(i_dcd_dec_2_init_mt_axi_s_awqos),
        .o_dcd_dec_2_init_mt_axi_s_awready(o_dcd_dec_2_init_mt_axi_s_awready),
        .i_dcd_dec_2_init_mt_axi_s_awsize(i_dcd_dec_2_init_mt_axi_s_awsize),
        .i_dcd_dec_2_init_mt_axi_s_awvalid(i_dcd_dec_2_init_mt_axi_s_awvalid),
        .o_dcd_dec_2_init_mt_axi_s_bid(o_dcd_dec_2_init_mt_axi_s_bid),
        .i_dcd_dec_2_init_mt_axi_s_bready(i_dcd_dec_2_init_mt_axi_s_bready),
        .o_dcd_dec_2_init_mt_axi_s_bresp(o_dcd_dec_2_init_mt_axi_s_bresp),
        .o_dcd_dec_2_init_mt_axi_s_bvalid(o_dcd_dec_2_init_mt_axi_s_bvalid),
        .i_dcd_dec_2_init_mt_axi_s_wdata(i_dcd_dec_2_init_mt_axi_s_wdata),
        .i_dcd_dec_2_init_mt_axi_s_wlast(i_dcd_dec_2_init_mt_axi_s_wlast),
        .o_dcd_dec_2_init_mt_axi_s_wready(o_dcd_dec_2_init_mt_axi_s_wready),
        .i_dcd_dec_2_init_mt_axi_s_wstrb(i_dcd_dec_2_init_mt_axi_s_wstrb),
        .i_dcd_dec_2_init_mt_axi_s_wvalid(i_dcd_dec_2_init_mt_axi_s_wvalid),
        .i_dcd_mcu_clk(i_dcd_mcu_clk),
        .i_dcd_mcu_clken(i_dcd_mcu_clken),
        .i_dcd_mcu_init_lt_axi_s_araddr(i_dcd_mcu_init_lt_axi_s_araddr),
        .i_dcd_mcu_init_lt_axi_s_arburst(i_dcd_mcu_init_lt_axi_s_arburst),
        .i_dcd_mcu_init_lt_axi_s_arcache(i_dcd_mcu_init_lt_axi_s_arcache),
        .i_dcd_mcu_init_lt_axi_s_arid(i_dcd_mcu_init_lt_axi_s_arid),
        .i_dcd_mcu_init_lt_axi_s_arlen(i_dcd_mcu_init_lt_axi_s_arlen),
        .i_dcd_mcu_init_lt_axi_s_arlock(i_dcd_mcu_init_lt_axi_s_arlock),
        .i_dcd_mcu_init_lt_axi_s_arprot(i_dcd_mcu_init_lt_axi_s_arprot),
        .i_dcd_mcu_init_lt_axi_s_arqos(i_dcd_mcu_init_lt_axi_s_arqos),
        .o_dcd_mcu_init_lt_axi_s_arready(o_dcd_mcu_init_lt_axi_s_arready),
        .i_dcd_mcu_init_lt_axi_s_arsize(i_dcd_mcu_init_lt_axi_s_arsize),
        .i_dcd_mcu_init_lt_axi_s_arvalid(i_dcd_mcu_init_lt_axi_s_arvalid),
        .o_dcd_mcu_init_lt_axi_s_rdata(o_dcd_mcu_init_lt_axi_s_rdata),
        .o_dcd_mcu_init_lt_axi_s_rid(o_dcd_mcu_init_lt_axi_s_rid),
        .o_dcd_mcu_init_lt_axi_s_rlast(o_dcd_mcu_init_lt_axi_s_rlast),
        .i_dcd_mcu_init_lt_axi_s_rready(i_dcd_mcu_init_lt_axi_s_rready),
        .o_dcd_mcu_init_lt_axi_s_rresp(o_dcd_mcu_init_lt_axi_s_rresp),
        .o_dcd_mcu_init_lt_axi_s_rvalid(o_dcd_mcu_init_lt_axi_s_rvalid),
        .i_dcd_mcu_init_lt_axi_s_awaddr(i_dcd_mcu_init_lt_axi_s_awaddr),
        .i_dcd_mcu_init_lt_axi_s_awburst(i_dcd_mcu_init_lt_axi_s_awburst),
        .i_dcd_mcu_init_lt_axi_s_awcache(i_dcd_mcu_init_lt_axi_s_awcache),
        .i_dcd_mcu_init_lt_axi_s_awid(i_dcd_mcu_init_lt_axi_s_awid),
        .i_dcd_mcu_init_lt_axi_s_awlen(i_dcd_mcu_init_lt_axi_s_awlen),
        .i_dcd_mcu_init_lt_axi_s_awlock(i_dcd_mcu_init_lt_axi_s_awlock),
        .i_dcd_mcu_init_lt_axi_s_awprot(i_dcd_mcu_init_lt_axi_s_awprot),
        .i_dcd_mcu_init_lt_axi_s_awqos(i_dcd_mcu_init_lt_axi_s_awqos),
        .o_dcd_mcu_init_lt_axi_s_awready(o_dcd_mcu_init_lt_axi_s_awready),
        .i_dcd_mcu_init_lt_axi_s_awsize(i_dcd_mcu_init_lt_axi_s_awsize),
        .i_dcd_mcu_init_lt_axi_s_awvalid(i_dcd_mcu_init_lt_axi_s_awvalid),
        .o_dcd_mcu_init_lt_axi_s_bid(o_dcd_mcu_init_lt_axi_s_bid),
        .i_dcd_mcu_init_lt_axi_s_bready(i_dcd_mcu_init_lt_axi_s_bready),
        .o_dcd_mcu_init_lt_axi_s_bresp(o_dcd_mcu_init_lt_axi_s_bresp),
        .o_dcd_mcu_init_lt_axi_s_bvalid(o_dcd_mcu_init_lt_axi_s_bvalid),
        .i_dcd_mcu_init_lt_axi_s_wdata(i_dcd_mcu_init_lt_axi_s_wdata),
        .i_dcd_mcu_init_lt_axi_s_wlast(i_dcd_mcu_init_lt_axi_s_wlast),
        .o_dcd_mcu_init_lt_axi_s_wready(o_dcd_mcu_init_lt_axi_s_wready),
        .i_dcd_mcu_init_lt_axi_s_wstrb(i_dcd_mcu_init_lt_axi_s_wstrb),
        .i_dcd_mcu_init_lt_axi_s_wvalid(i_dcd_mcu_init_lt_axi_s_wvalid),
        .o_dcd_mcu_pwr_idle_val(o_dcd_mcu_pwr_idle_val),
        .o_dcd_mcu_pwr_idle_ack(o_dcd_mcu_pwr_idle_ack),
        .i_dcd_mcu_pwr_idle_req(i_dcd_mcu_pwr_idle_req),
        .i_dcd_mcu_rst_n(i_dcd_mcu_rst_n),
        .o_dcd_pwr_idle_val(o_dcd_pwr_idle_val),
        .o_dcd_pwr_idle_ack(o_dcd_pwr_idle_ack),
        .i_dcd_pwr_idle_req(i_dcd_pwr_idle_req),
        .o_dcd_targ_cfg_apb_m_paddr(o_dcd_targ_cfg_apb_m_paddr),
        .o_dcd_targ_cfg_apb_m_penable(o_dcd_targ_cfg_apb_m_penable),
        .o_dcd_targ_cfg_apb_m_pprot(o_dcd_targ_cfg_apb_m_pprot),
        .i_dcd_targ_cfg_apb_m_prdata(i_dcd_targ_cfg_apb_m_prdata),
        .i_dcd_targ_cfg_apb_m_pready(i_dcd_targ_cfg_apb_m_pready),
        .o_dcd_targ_cfg_apb_m_psel(o_dcd_targ_cfg_apb_m_psel),
        .i_dcd_targ_cfg_apb_m_pslverr(i_dcd_targ_cfg_apb_m_pslverr),
        .o_dcd_targ_cfg_apb_m_pstrb(o_dcd_targ_cfg_apb_m_pstrb),
        .o_dcd_targ_cfg_apb_m_pwdata(o_dcd_targ_cfg_apb_m_pwdata),
        .o_dcd_targ_cfg_apb_m_pwrite(o_dcd_targ_cfg_apb_m_pwrite),
        .o_dcd_targ_syscfg_apb_m_paddr(o_dcd_targ_syscfg_apb_m_paddr),
        .o_dcd_targ_syscfg_apb_m_penable(o_dcd_targ_syscfg_apb_m_penable),
        .o_dcd_targ_syscfg_apb_m_pprot(o_dcd_targ_syscfg_apb_m_pprot),
        .i_dcd_targ_syscfg_apb_m_prdata(i_dcd_targ_syscfg_apb_m_prdata),
        .i_dcd_targ_syscfg_apb_m_pready(i_dcd_targ_syscfg_apb_m_pready),
        .o_dcd_targ_syscfg_apb_m_psel(o_dcd_targ_syscfg_apb_m_psel),
        .i_dcd_targ_syscfg_apb_m_pslverr(i_dcd_targ_syscfg_apb_m_pslverr),
        .o_dcd_targ_syscfg_apb_m_pstrb(o_dcd_targ_syscfg_apb_m_pstrb),
        .o_dcd_targ_syscfg_apb_m_pwdata(o_dcd_targ_syscfg_apb_m_pwdata),
        .o_dcd_targ_syscfg_apb_m_pwrite(o_dcd_targ_syscfg_apb_m_pwrite),
        .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_data),
        .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_head),
        .o_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_rdy),
        .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_tail),
        .i_dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld(dp_lnk_cross_east_to_soc_512_0_egr_wr_req_to_lnk_cross_east_to_soc_512_0_ingr_wr_req_vld),
        .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_data),
        .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_head),
        .i_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld(dp_lnk_cross_east_to_soc_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_0_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_data),
        .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_head),
        .o_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_rdy),
        .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_tail),
        .i_dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld(dp_lnk_cross_east_to_soc_512_1_egr_wr_req_to_lnk_cross_east_to_soc_512_1_ingr_wr_req_vld),
        .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_data),
        .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_head),
        .i_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld(dp_lnk_cross_east_to_soc_512_1_ingr_wr_req_resp_to_lnk_cross_east_to_soc_512_1_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_data),
        .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_head),
        .o_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_rdy),
        .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_tail),
        .i_dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld(dp_lnk_cross_east_to_soc_512_2_egr_rd_req_to_lnk_cross_east_to_soc_512_2_ingr_rd_req_vld),
        .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_data),
        .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_head),
        .i_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld(dp_lnk_cross_east_to_soc_512_2_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_2_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_data),
        .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_head),
        .o_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_rdy),
        .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_tail),
        .i_dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld(dp_lnk_cross_east_to_soc_512_3_egr_rd_req_to_lnk_cross_east_to_soc_512_3_ingr_rd_req_vld),
        .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_data),
        .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_head),
        .i_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld(dp_lnk_cross_east_to_soc_512_3_ingr_rd_req_resp_to_lnk_cross_east_to_soc_512_3_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_data),
        .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_head),
        .o_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_rdy),
        .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_tail),
        .i_dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld(dp_lnk_cross_east_to_soc_64_egr_req_to_lnk_cross_east_to_soc_64_ingr_req_vld),
        .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_data),
        .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_head),
        .i_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_tail),
        .o_dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld(dp_lnk_cross_east_to_soc_64_ingr_req_resp_to_lnk_cross_east_to_soc_64_egr_req_resp_vld),
        .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_data),
        .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_head),
        .o_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_rdy),
        .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_tail),
        .i_dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld(dp_lnk_cross_soc_periph_to_soc_64_egr_to_lnk_cross_soc_periph_to_soc_64_ingr_req_vld),
        .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_data),
        .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_head),
        .i_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_rdy),
        .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_tail),
        .o_dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld(dp_lnk_cross_soc_periph_to_soc_64_ingr_req_resp_to_lnk_cross_soc_periph_to_soc_64_egr_resp_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_data),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_head),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_256_0_egr_req_to_lnk_cross_soc_to_ddr_e_256_0_ingr_req_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_data),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_head),
        .o_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_256_0_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_0_egr_req_resp_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_data),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_head),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_256_1_egr_req_to_lnk_cross_soc_to_ddr_e_256_1_ingr_req_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_data),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_head),
        .o_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_256_1_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_1_egr_req_resp_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_data),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_head),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_256_2_egr_req_to_lnk_cross_soc_to_ddr_e_256_2_ingr_req_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_data),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_head),
        .o_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_256_2_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_2_egr_req_resp_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_data),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_head),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_256_3_egr_req_to_lnk_cross_soc_to_ddr_e_256_3_ingr_req_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_data),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_head),
        .o_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_256_3_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_256_3_egr_req_resp_vld),
        .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_data),
        .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_head),
        .i_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_rdy),
        .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_tail),
        .o_dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld(dp_lnk_cross_soc_to_ddr_e_64_egr_req_to_lnk_cross_soc_to_ddr_e_64_ingr_req_vld),
        .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_data),
        .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_head),
        .o_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_tail),
        .i_dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld(dp_lnk_cross_soc_to_ddr_e_64_ingr_req_resp_to_lnk_cross_soc_to_ddr_e_64_egr_req_resp_vld),
        .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_data),
        .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_head),
        .i_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_rdy),
        .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_tail),
        .o_dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld(dp_lnk_cross_soc_to_east_512_0_egr_wr_req_to_lnk_cross_soc_to_east_512_0_ingr_wr_req_vld),
        .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_data),
        .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_head),
        .o_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld(dp_lnk_cross_soc_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_soc_to_east_512_0_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_data),
        .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_head),
        .i_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_rdy),
        .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_tail),
        .o_dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld(dp_lnk_cross_soc_to_east_512_1_egr_rd_req_to_lnk_cross_soc_to_east_512_1_ingr_rd_req_vld),
        .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_data),
        .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_head),
        .o_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld(dp_lnk_cross_soc_to_east_512_1_ingr_rd_req_resp_to_lnk_cross_soc_to_east_512_1_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_data),
        .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_head),
        .i_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_rdy),
        .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_tail),
        .o_dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld(dp_lnk_cross_soc_to_east_64_egr_req_to_lnk_cross_soc_to_east_64_ingr_req_vld),
        .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_data),
        .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_head),
        .o_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_tail),
        .i_dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld(dp_lnk_cross_soc_to_east_64_ingr_req_resp_to_lnk_cross_soc_to_east_64_egr_req_resp_vld),
        .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
        .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
        .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
        .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
        .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
        .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
        .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
        .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
        .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
        .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
        .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
        .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),
        .i_noc_clk(i_noc_clk),
        .i_noc_rst_n(i_noc_rst_n),
        .i_pcie_aon_clk(i_pcie_aon_clk),
        .i_pcie_aon_rst_n(i_pcie_aon_rst_n),
        .i_pcie_init_mt_clk(i_pcie_init_mt_clk),
        .i_pcie_init_mt_clken(i_pcie_init_mt_clken),
        .o_pcie_init_mt_pwr_idle_val(o_pcie_init_mt_pwr_idle_val),
        .o_pcie_init_mt_pwr_idle_ack(o_pcie_init_mt_pwr_idle_ack),
        .i_pcie_init_mt_pwr_idle_req(i_pcie_init_mt_pwr_idle_req),
        .i_pcie_init_mt_axi_s_araddr(i_pcie_init_mt_axi_s_araddr),
        .i_pcie_init_mt_axi_s_arburst(i_pcie_init_mt_axi_s_arburst),
        .i_pcie_init_mt_axi_s_arcache(i_pcie_init_mt_axi_s_arcache),
        .i_pcie_init_mt_axi_s_arid(i_pcie_init_mt_axi_s_arid),
        .i_pcie_init_mt_axi_s_arlen(i_pcie_init_mt_axi_s_arlen),
        .i_pcie_init_mt_axi_s_arlock(i_pcie_init_mt_axi_s_arlock),
        .i_pcie_init_mt_axi_s_arprot(i_pcie_init_mt_axi_s_arprot),
        .i_pcie_init_mt_axi_s_arqos(i_pcie_init_mt_axi_s_arqos),
        .o_pcie_init_mt_axi_s_arready(o_pcie_init_mt_axi_s_arready),
        .i_pcie_init_mt_axi_s_arsize(i_pcie_init_mt_axi_s_arsize),
        .i_pcie_init_mt_axi_s_arvalid(i_pcie_init_mt_axi_s_arvalid),
        .o_pcie_init_mt_axi_s_rdata(o_pcie_init_mt_axi_s_rdata),
        .o_pcie_init_mt_axi_s_rid(o_pcie_init_mt_axi_s_rid),
        .o_pcie_init_mt_axi_s_rlast(o_pcie_init_mt_axi_s_rlast),
        .i_pcie_init_mt_axi_s_rready(i_pcie_init_mt_axi_s_rready),
        .o_pcie_init_mt_axi_s_rresp(o_pcie_init_mt_axi_s_rresp),
        .o_pcie_init_mt_axi_s_rvalid(o_pcie_init_mt_axi_s_rvalid),
        .i_pcie_init_mt_rst_n(i_pcie_init_mt_rst_n),
        .i_pcie_init_mt_axi_s_awaddr(i_pcie_init_mt_axi_s_awaddr),
        .i_pcie_init_mt_axi_s_awburst(i_pcie_init_mt_axi_s_awburst),
        .i_pcie_init_mt_axi_s_awcache(i_pcie_init_mt_axi_s_awcache),
        .i_pcie_init_mt_axi_s_awid(i_pcie_init_mt_axi_s_awid),
        .i_pcie_init_mt_axi_s_awlen(i_pcie_init_mt_axi_s_awlen),
        .i_pcie_init_mt_axi_s_awlock(i_pcie_init_mt_axi_s_awlock),
        .i_pcie_init_mt_axi_s_awprot(i_pcie_init_mt_axi_s_awprot),
        .i_pcie_init_mt_axi_s_awqos(i_pcie_init_mt_axi_s_awqos),
        .o_pcie_init_mt_axi_s_awready(o_pcie_init_mt_axi_s_awready),
        .i_pcie_init_mt_axi_s_awsize(i_pcie_init_mt_axi_s_awsize),
        .i_pcie_init_mt_axi_s_awvalid(i_pcie_init_mt_axi_s_awvalid),
        .o_pcie_init_mt_axi_s_bid(o_pcie_init_mt_axi_s_bid),
        .i_pcie_init_mt_axi_s_bready(i_pcie_init_mt_axi_s_bready),
        .o_pcie_init_mt_axi_s_bresp(o_pcie_init_mt_axi_s_bresp),
        .o_pcie_init_mt_axi_s_bvalid(o_pcie_init_mt_axi_s_bvalid),
        .i_pcie_init_mt_axi_s_wdata(i_pcie_init_mt_axi_s_wdata),
        .i_pcie_init_mt_axi_s_wlast(i_pcie_init_mt_axi_s_wlast),
        .o_pcie_init_mt_axi_s_wready(o_pcie_init_mt_axi_s_wready),
        .i_pcie_init_mt_axi_s_wstrb(i_pcie_init_mt_axi_s_wstrb),
        .i_pcie_init_mt_axi_s_wvalid(i_pcie_init_mt_axi_s_wvalid),
        .o_pcie_targ_cfg_apb_m_paddr(o_pcie_targ_cfg_apb_m_paddr),
        .o_pcie_targ_cfg_apb_m_penable(o_pcie_targ_cfg_apb_m_penable),
        .o_pcie_targ_cfg_apb_m_pprot(o_pcie_targ_cfg_apb_m_pprot),
        .i_pcie_targ_cfg_apb_m_prdata(i_pcie_targ_cfg_apb_m_prdata),
        .i_pcie_targ_cfg_apb_m_pready(i_pcie_targ_cfg_apb_m_pready),
        .o_pcie_targ_cfg_apb_m_psel(o_pcie_targ_cfg_apb_m_psel),
        .i_pcie_targ_cfg_apb_m_pslverr(i_pcie_targ_cfg_apb_m_pslverr),
        .o_pcie_targ_cfg_apb_m_pstrb(o_pcie_targ_cfg_apb_m_pstrb),
        .o_pcie_targ_cfg_apb_m_pwdata(o_pcie_targ_cfg_apb_m_pwdata),
        .o_pcie_targ_cfg_apb_m_pwrite(o_pcie_targ_cfg_apb_m_pwrite),
        .i_pcie_targ_cfg_clk(i_pcie_targ_cfg_clk),
        .i_pcie_targ_cfg_clken(i_pcie_targ_cfg_clken),
        .o_pcie_targ_cfg_dbi_axi_m_araddr(o_pcie_targ_cfg_dbi_axi_m_araddr),
        .o_pcie_targ_cfg_dbi_axi_m_arburst(o_pcie_targ_cfg_dbi_axi_m_arburst),
        .o_pcie_targ_cfg_dbi_axi_m_arcache(o_pcie_targ_cfg_dbi_axi_m_arcache),
        .o_pcie_targ_cfg_dbi_axi_m_arid(o_pcie_targ_cfg_dbi_axi_m_arid),
        .o_pcie_targ_cfg_dbi_axi_m_arlen(o_pcie_targ_cfg_dbi_axi_m_arlen),
        .o_pcie_targ_cfg_dbi_axi_m_arlock(o_pcie_targ_cfg_dbi_axi_m_arlock),
        .o_pcie_targ_cfg_dbi_axi_m_arprot(o_pcie_targ_cfg_dbi_axi_m_arprot),
        .o_pcie_targ_cfg_dbi_axi_m_arqos(o_pcie_targ_cfg_dbi_axi_m_arqos),
        .i_pcie_targ_cfg_dbi_axi_m_arready(i_pcie_targ_cfg_dbi_axi_m_arready),
        .o_pcie_targ_cfg_dbi_axi_m_arsize(o_pcie_targ_cfg_dbi_axi_m_arsize),
        .o_pcie_targ_cfg_dbi_axi_m_arvalid(o_pcie_targ_cfg_dbi_axi_m_arvalid),
        .o_pcie_targ_cfg_dbi_axi_m_awaddr(o_pcie_targ_cfg_dbi_axi_m_awaddr),
        .o_pcie_targ_cfg_dbi_axi_m_awburst(o_pcie_targ_cfg_dbi_axi_m_awburst),
        .o_pcie_targ_cfg_dbi_axi_m_awcache(o_pcie_targ_cfg_dbi_axi_m_awcache),
        .o_pcie_targ_cfg_dbi_axi_m_awid(o_pcie_targ_cfg_dbi_axi_m_awid),
        .o_pcie_targ_cfg_dbi_axi_m_awlen(o_pcie_targ_cfg_dbi_axi_m_awlen),
        .o_pcie_targ_cfg_dbi_axi_m_awlock(o_pcie_targ_cfg_dbi_axi_m_awlock),
        .o_pcie_targ_cfg_dbi_axi_m_awprot(o_pcie_targ_cfg_dbi_axi_m_awprot),
        .o_pcie_targ_cfg_dbi_axi_m_awqos(o_pcie_targ_cfg_dbi_axi_m_awqos),
        .i_pcie_targ_cfg_dbi_axi_m_awready(i_pcie_targ_cfg_dbi_axi_m_awready),
        .o_pcie_targ_cfg_dbi_axi_m_awsize(o_pcie_targ_cfg_dbi_axi_m_awsize),
        .o_pcie_targ_cfg_dbi_axi_m_awvalid(o_pcie_targ_cfg_dbi_axi_m_awvalid),
        .i_pcie_targ_cfg_dbi_axi_m_bid(i_pcie_targ_cfg_dbi_axi_m_bid),
        .o_pcie_targ_cfg_dbi_axi_m_bready(o_pcie_targ_cfg_dbi_axi_m_bready),
        .i_pcie_targ_cfg_dbi_axi_m_bresp(i_pcie_targ_cfg_dbi_axi_m_bresp),
        .i_pcie_targ_cfg_dbi_axi_m_bvalid(i_pcie_targ_cfg_dbi_axi_m_bvalid),
        .i_pcie_targ_cfg_dbi_axi_m_rdata(i_pcie_targ_cfg_dbi_axi_m_rdata),
        .i_pcie_targ_cfg_dbi_axi_m_rid(i_pcie_targ_cfg_dbi_axi_m_rid),
        .i_pcie_targ_cfg_dbi_axi_m_rlast(i_pcie_targ_cfg_dbi_axi_m_rlast),
        .o_pcie_targ_cfg_dbi_axi_m_rready(o_pcie_targ_cfg_dbi_axi_m_rready),
        .i_pcie_targ_cfg_dbi_axi_m_rresp(i_pcie_targ_cfg_dbi_axi_m_rresp),
        .i_pcie_targ_cfg_dbi_axi_m_rvalid(i_pcie_targ_cfg_dbi_axi_m_rvalid),
        .o_pcie_targ_cfg_dbi_axi_m_wdata(o_pcie_targ_cfg_dbi_axi_m_wdata),
        .o_pcie_targ_cfg_dbi_axi_m_wlast(o_pcie_targ_cfg_dbi_axi_m_wlast),
        .i_pcie_targ_cfg_dbi_axi_m_wready(i_pcie_targ_cfg_dbi_axi_m_wready),
        .o_pcie_targ_cfg_dbi_axi_m_wstrb(o_pcie_targ_cfg_dbi_axi_m_wstrb),
        .o_pcie_targ_cfg_dbi_axi_m_wvalid(o_pcie_targ_cfg_dbi_axi_m_wvalid),
        .i_pcie_targ_cfg_dbi_clk(i_pcie_targ_cfg_dbi_clk),
        .i_pcie_targ_cfg_dbi_clken(i_pcie_targ_cfg_dbi_clken),
        .o_pcie_targ_cfg_dbi_pwr_idle_val(o_pcie_targ_cfg_dbi_pwr_idle_val),
        .o_pcie_targ_cfg_dbi_pwr_idle_ack(o_pcie_targ_cfg_dbi_pwr_idle_ack),
        .i_pcie_targ_cfg_dbi_pwr_idle_req(i_pcie_targ_cfg_dbi_pwr_idle_req),
        .i_pcie_targ_cfg_dbi_rst_n(i_pcie_targ_cfg_dbi_rst_n),
        .o_pcie_targ_cfg_pwr_idle_val(o_pcie_targ_cfg_pwr_idle_val),
        .o_pcie_targ_cfg_pwr_idle_ack(o_pcie_targ_cfg_pwr_idle_ack),
        .i_pcie_targ_cfg_pwr_idle_req(i_pcie_targ_cfg_pwr_idle_req),
        .i_pcie_targ_cfg_rst_n(i_pcie_targ_cfg_rst_n),
        .i_pcie_targ_mt_clk(i_pcie_targ_mt_clk),
        .i_pcie_targ_mt_clken(i_pcie_targ_mt_clken),
        .o_pcie_targ_mt_pwr_idle_val(o_pcie_targ_mt_pwr_idle_val),
        .o_pcie_targ_mt_pwr_idle_ack(o_pcie_targ_mt_pwr_idle_ack),
        .i_pcie_targ_mt_pwr_idle_req(i_pcie_targ_mt_pwr_idle_req),
        .o_pcie_targ_mt_axi_m_araddr(o_pcie_targ_mt_axi_m_araddr),
        .o_pcie_targ_mt_axi_m_arburst(o_pcie_targ_mt_axi_m_arburst),
        .o_pcie_targ_mt_axi_m_arcache(o_pcie_targ_mt_axi_m_arcache),
        .o_pcie_targ_mt_axi_m_arid(o_pcie_targ_mt_axi_m_arid),
        .o_pcie_targ_mt_axi_m_arlen(o_pcie_targ_mt_axi_m_arlen),
        .o_pcie_targ_mt_axi_m_arlock(o_pcie_targ_mt_axi_m_arlock),
        .o_pcie_targ_mt_axi_m_arprot(o_pcie_targ_mt_axi_m_arprot),
        .o_pcie_targ_mt_axi_m_arqos(o_pcie_targ_mt_axi_m_arqos),
        .i_pcie_targ_mt_axi_m_arready(i_pcie_targ_mt_axi_m_arready),
        .o_pcie_targ_mt_axi_m_arsize(o_pcie_targ_mt_axi_m_arsize),
        .o_pcie_targ_mt_axi_m_arvalid(o_pcie_targ_mt_axi_m_arvalid),
        .i_pcie_targ_mt_axi_m_rdata(i_pcie_targ_mt_axi_m_rdata),
        .i_pcie_targ_mt_axi_m_rid(i_pcie_targ_mt_axi_m_rid),
        .i_pcie_targ_mt_axi_m_rlast(i_pcie_targ_mt_axi_m_rlast),
        .o_pcie_targ_mt_axi_m_rready(o_pcie_targ_mt_axi_m_rready),
        .i_pcie_targ_mt_axi_m_rresp(i_pcie_targ_mt_axi_m_rresp),
        .i_pcie_targ_mt_axi_m_rvalid(i_pcie_targ_mt_axi_m_rvalid),
        .i_pcie_targ_mt_rst_n(i_pcie_targ_mt_rst_n),
        .o_pcie_targ_mt_axi_m_awaddr(o_pcie_targ_mt_axi_m_awaddr),
        .o_pcie_targ_mt_axi_m_awburst(o_pcie_targ_mt_axi_m_awburst),
        .o_pcie_targ_mt_axi_m_awcache(o_pcie_targ_mt_axi_m_awcache),
        .o_pcie_targ_mt_axi_m_awid(o_pcie_targ_mt_axi_m_awid),
        .o_pcie_targ_mt_axi_m_awlen(o_pcie_targ_mt_axi_m_awlen),
        .o_pcie_targ_mt_axi_m_awlock(o_pcie_targ_mt_axi_m_awlock),
        .o_pcie_targ_mt_axi_m_awprot(o_pcie_targ_mt_axi_m_awprot),
        .o_pcie_targ_mt_axi_m_awqos(o_pcie_targ_mt_axi_m_awqos),
        .i_pcie_targ_mt_axi_m_awready(i_pcie_targ_mt_axi_m_awready),
        .o_pcie_targ_mt_axi_m_awsize(o_pcie_targ_mt_axi_m_awsize),
        .o_pcie_targ_mt_axi_m_awvalid(o_pcie_targ_mt_axi_m_awvalid),
        .i_pcie_targ_mt_axi_m_bid(i_pcie_targ_mt_axi_m_bid),
        .o_pcie_targ_mt_axi_m_bready(o_pcie_targ_mt_axi_m_bready),
        .i_pcie_targ_mt_axi_m_bresp(i_pcie_targ_mt_axi_m_bresp),
        .i_pcie_targ_mt_axi_m_bvalid(i_pcie_targ_mt_axi_m_bvalid),
        .o_pcie_targ_mt_axi_m_wdata(o_pcie_targ_mt_axi_m_wdata),
        .o_pcie_targ_mt_axi_m_wlast(o_pcie_targ_mt_axi_m_wlast),
        .i_pcie_targ_mt_axi_m_wready(i_pcie_targ_mt_axi_m_wready),
        .o_pcie_targ_mt_axi_m_wstrb(o_pcie_targ_mt_axi_m_wstrb),
        .o_pcie_targ_mt_axi_m_wvalid(o_pcie_targ_mt_axi_m_wvalid),
        .o_pcie_targ_syscfg_apb_m_paddr(o_pcie_targ_syscfg_apb_m_paddr),
        .o_pcie_targ_syscfg_apb_m_penable(o_pcie_targ_syscfg_apb_m_penable),
        .o_pcie_targ_syscfg_apb_m_pprot(o_pcie_targ_syscfg_apb_m_pprot),
        .i_pcie_targ_syscfg_apb_m_prdata(i_pcie_targ_syscfg_apb_m_prdata),
        .i_pcie_targ_syscfg_apb_m_pready(i_pcie_targ_syscfg_apb_m_pready),
        .o_pcie_targ_syscfg_apb_m_psel(o_pcie_targ_syscfg_apb_m_psel),
        .i_pcie_targ_syscfg_apb_m_pslverr(i_pcie_targ_syscfg_apb_m_pslverr),
        .o_pcie_targ_syscfg_apb_m_pstrb(o_pcie_targ_syscfg_apb_m_pstrb),
        .o_pcie_targ_syscfg_apb_m_pwdata(o_pcie_targ_syscfg_apb_m_pwdata),
        .o_pcie_targ_syscfg_apb_m_pwrite(o_pcie_targ_syscfg_apb_m_pwrite),
        .i_pve_0_aon_clk(i_pve_0_aon_clk),
        .i_pve_0_aon_rst_n(i_pve_0_aon_rst_n),
        .i_pve_0_clk(i_pve_0_clk),
        .i_pve_0_clken(i_pve_0_clken),
        .i_pve_0_init_ht_axi_s_araddr(i_pve_0_init_ht_axi_s_araddr),
        .i_pve_0_init_ht_axi_s_arburst(i_pve_0_init_ht_axi_s_arburst),
        .i_pve_0_init_ht_axi_s_arcache(i_pve_0_init_ht_axi_s_arcache),
        .i_pve_0_init_ht_axi_s_arid(i_pve_0_init_ht_axi_s_arid),
        .i_pve_0_init_ht_axi_s_arlen(i_pve_0_init_ht_axi_s_arlen),
        .i_pve_0_init_ht_axi_s_arlock(i_pve_0_init_ht_axi_s_arlock),
        .i_pve_0_init_ht_axi_s_arprot(i_pve_0_init_ht_axi_s_arprot),
        .o_pve_0_init_ht_axi_s_arready(o_pve_0_init_ht_axi_s_arready),
        .i_pve_0_init_ht_axi_s_arsize(i_pve_0_init_ht_axi_s_arsize),
        .i_pve_0_init_ht_axi_s_arvalid(i_pve_0_init_ht_axi_s_arvalid),
        .o_pve_0_init_ht_axi_s_rdata(o_pve_0_init_ht_axi_s_rdata),
        .o_pve_0_init_ht_axi_s_rid(o_pve_0_init_ht_axi_s_rid),
        .o_pve_0_init_ht_axi_s_rlast(o_pve_0_init_ht_axi_s_rlast),
        .i_pve_0_init_ht_axi_s_rready(i_pve_0_init_ht_axi_s_rready),
        .o_pve_0_init_ht_axi_s_rresp(o_pve_0_init_ht_axi_s_rresp),
        .o_pve_0_init_ht_axi_s_rvalid(o_pve_0_init_ht_axi_s_rvalid),
        .i_pve_0_init_ht_axi_s_awaddr(i_pve_0_init_ht_axi_s_awaddr),
        .i_pve_0_init_ht_axi_s_awburst(i_pve_0_init_ht_axi_s_awburst),
        .i_pve_0_init_ht_axi_s_awcache(i_pve_0_init_ht_axi_s_awcache),
        .i_pve_0_init_ht_axi_s_awid(i_pve_0_init_ht_axi_s_awid),
        .i_pve_0_init_ht_axi_s_awlen(i_pve_0_init_ht_axi_s_awlen),
        .i_pve_0_init_ht_axi_s_awlock(i_pve_0_init_ht_axi_s_awlock),
        .i_pve_0_init_ht_axi_s_awprot(i_pve_0_init_ht_axi_s_awprot),
        .o_pve_0_init_ht_axi_s_awready(o_pve_0_init_ht_axi_s_awready),
        .i_pve_0_init_ht_axi_s_awsize(i_pve_0_init_ht_axi_s_awsize),
        .i_pve_0_init_ht_axi_s_awvalid(i_pve_0_init_ht_axi_s_awvalid),
        .o_pve_0_init_ht_axi_s_bid(o_pve_0_init_ht_axi_s_bid),
        .i_pve_0_init_ht_axi_s_bready(i_pve_0_init_ht_axi_s_bready),
        .o_pve_0_init_ht_axi_s_bresp(o_pve_0_init_ht_axi_s_bresp),
        .o_pve_0_init_ht_axi_s_bvalid(o_pve_0_init_ht_axi_s_bvalid),
        .i_pve_0_init_ht_axi_s_wdata(i_pve_0_init_ht_axi_s_wdata),
        .i_pve_0_init_ht_axi_s_wlast(i_pve_0_init_ht_axi_s_wlast),
        .o_pve_0_init_ht_axi_s_wready(o_pve_0_init_ht_axi_s_wready),
        .i_pve_0_init_ht_axi_s_wstrb(i_pve_0_init_ht_axi_s_wstrb),
        .i_pve_0_init_ht_axi_s_wvalid(i_pve_0_init_ht_axi_s_wvalid),
        .i_pve_0_init_lt_axi_s_araddr(i_pve_0_init_lt_axi_s_araddr),
        .i_pve_0_init_lt_axi_s_arburst(i_pve_0_init_lt_axi_s_arburst),
        .i_pve_0_init_lt_axi_s_arcache(i_pve_0_init_lt_axi_s_arcache),
        .i_pve_0_init_lt_axi_s_arid(i_pve_0_init_lt_axi_s_arid),
        .i_pve_0_init_lt_axi_s_arlen(i_pve_0_init_lt_axi_s_arlen),
        .i_pve_0_init_lt_axi_s_arlock(i_pve_0_init_lt_axi_s_arlock),
        .i_pve_0_init_lt_axi_s_arprot(i_pve_0_init_lt_axi_s_arprot),
        .i_pve_0_init_lt_axi_s_arqos(i_pve_0_init_lt_axi_s_arqos),
        .o_pve_0_init_lt_axi_s_arready(o_pve_0_init_lt_axi_s_arready),
        .i_pve_0_init_lt_axi_s_arsize(i_pve_0_init_lt_axi_s_arsize),
        .i_pve_0_init_lt_axi_s_arvalid(i_pve_0_init_lt_axi_s_arvalid),
        .o_pve_0_init_lt_axi_s_rdata(o_pve_0_init_lt_axi_s_rdata),
        .o_pve_0_init_lt_axi_s_rid(o_pve_0_init_lt_axi_s_rid),
        .o_pve_0_init_lt_axi_s_rlast(o_pve_0_init_lt_axi_s_rlast),
        .i_pve_0_init_lt_axi_s_rready(i_pve_0_init_lt_axi_s_rready),
        .o_pve_0_init_lt_axi_s_rresp(o_pve_0_init_lt_axi_s_rresp),
        .o_pve_0_init_lt_axi_s_rvalid(o_pve_0_init_lt_axi_s_rvalid),
        .i_pve_0_init_lt_axi_s_awaddr(i_pve_0_init_lt_axi_s_awaddr),
        .i_pve_0_init_lt_axi_s_awburst(i_pve_0_init_lt_axi_s_awburst),
        .i_pve_0_init_lt_axi_s_awcache(i_pve_0_init_lt_axi_s_awcache),
        .i_pve_0_init_lt_axi_s_awid(i_pve_0_init_lt_axi_s_awid),
        .i_pve_0_init_lt_axi_s_awlen(i_pve_0_init_lt_axi_s_awlen),
        .i_pve_0_init_lt_axi_s_awlock(i_pve_0_init_lt_axi_s_awlock),
        .i_pve_0_init_lt_axi_s_awprot(i_pve_0_init_lt_axi_s_awprot),
        .i_pve_0_init_lt_axi_s_awqos(i_pve_0_init_lt_axi_s_awqos),
        .o_pve_0_init_lt_axi_s_awready(o_pve_0_init_lt_axi_s_awready),
        .i_pve_0_init_lt_axi_s_awsize(i_pve_0_init_lt_axi_s_awsize),
        .i_pve_0_init_lt_axi_s_awvalid(i_pve_0_init_lt_axi_s_awvalid),
        .o_pve_0_init_lt_axi_s_bid(o_pve_0_init_lt_axi_s_bid),
        .i_pve_0_init_lt_axi_s_bready(i_pve_0_init_lt_axi_s_bready),
        .o_pve_0_init_lt_axi_s_bresp(o_pve_0_init_lt_axi_s_bresp),
        .o_pve_0_init_lt_axi_s_bvalid(o_pve_0_init_lt_axi_s_bvalid),
        .i_pve_0_init_lt_axi_s_wdata(i_pve_0_init_lt_axi_s_wdata),
        .i_pve_0_init_lt_axi_s_wlast(i_pve_0_init_lt_axi_s_wlast),
        .o_pve_0_init_lt_axi_s_wready(o_pve_0_init_lt_axi_s_wready),
        .i_pve_0_init_lt_axi_s_wstrb(i_pve_0_init_lt_axi_s_wstrb),
        .i_pve_0_init_lt_axi_s_wvalid(i_pve_0_init_lt_axi_s_wvalid),
        .o_pve_0_pwr_idle_val(o_pve_0_pwr_idle_val),
        .o_pve_0_pwr_idle_ack(o_pve_0_pwr_idle_ack),
        .i_pve_0_pwr_idle_req(i_pve_0_pwr_idle_req),
        .i_pve_0_rst_n(i_pve_0_rst_n),
        .o_pve_0_targ_lt_axi_m_araddr(o_pve_0_targ_lt_axi_m_araddr),
        .o_pve_0_targ_lt_axi_m_arburst(o_pve_0_targ_lt_axi_m_arburst),
        .o_pve_0_targ_lt_axi_m_arcache(o_pve_0_targ_lt_axi_m_arcache),
        .o_pve_0_targ_lt_axi_m_arid(o_pve_0_targ_lt_axi_m_arid),
        .o_pve_0_targ_lt_axi_m_arlen(o_pve_0_targ_lt_axi_m_arlen),
        .o_pve_0_targ_lt_axi_m_arlock(o_pve_0_targ_lt_axi_m_arlock),
        .o_pve_0_targ_lt_axi_m_arprot(o_pve_0_targ_lt_axi_m_arprot),
        .o_pve_0_targ_lt_axi_m_arqos(o_pve_0_targ_lt_axi_m_arqos),
        .i_pve_0_targ_lt_axi_m_arready(i_pve_0_targ_lt_axi_m_arready),
        .o_pve_0_targ_lt_axi_m_arsize(o_pve_0_targ_lt_axi_m_arsize),
        .o_pve_0_targ_lt_axi_m_arvalid(o_pve_0_targ_lt_axi_m_arvalid),
        .o_pve_0_targ_lt_axi_m_awaddr(o_pve_0_targ_lt_axi_m_awaddr),
        .o_pve_0_targ_lt_axi_m_awburst(o_pve_0_targ_lt_axi_m_awburst),
        .o_pve_0_targ_lt_axi_m_awcache(o_pve_0_targ_lt_axi_m_awcache),
        .o_pve_0_targ_lt_axi_m_awid(o_pve_0_targ_lt_axi_m_awid),
        .o_pve_0_targ_lt_axi_m_awlen(o_pve_0_targ_lt_axi_m_awlen),
        .o_pve_0_targ_lt_axi_m_awlock(o_pve_0_targ_lt_axi_m_awlock),
        .o_pve_0_targ_lt_axi_m_awprot(o_pve_0_targ_lt_axi_m_awprot),
        .o_pve_0_targ_lt_axi_m_awqos(o_pve_0_targ_lt_axi_m_awqos),
        .i_pve_0_targ_lt_axi_m_awready(i_pve_0_targ_lt_axi_m_awready),
        .o_pve_0_targ_lt_axi_m_awsize(o_pve_0_targ_lt_axi_m_awsize),
        .o_pve_0_targ_lt_axi_m_awvalid(o_pve_0_targ_lt_axi_m_awvalid),
        .i_pve_0_targ_lt_axi_m_bid(i_pve_0_targ_lt_axi_m_bid),
        .o_pve_0_targ_lt_axi_m_bready(o_pve_0_targ_lt_axi_m_bready),
        .i_pve_0_targ_lt_axi_m_bresp(i_pve_0_targ_lt_axi_m_bresp),
        .i_pve_0_targ_lt_axi_m_bvalid(i_pve_0_targ_lt_axi_m_bvalid),
        .i_pve_0_targ_lt_axi_m_rdata(i_pve_0_targ_lt_axi_m_rdata),
        .i_pve_0_targ_lt_axi_m_rid(i_pve_0_targ_lt_axi_m_rid),
        .i_pve_0_targ_lt_axi_m_rlast(i_pve_0_targ_lt_axi_m_rlast),
        .o_pve_0_targ_lt_axi_m_rready(o_pve_0_targ_lt_axi_m_rready),
        .i_pve_0_targ_lt_axi_m_rresp(i_pve_0_targ_lt_axi_m_rresp),
        .i_pve_0_targ_lt_axi_m_rvalid(i_pve_0_targ_lt_axi_m_rvalid),
        .o_pve_0_targ_lt_axi_m_wdata(o_pve_0_targ_lt_axi_m_wdata),
        .o_pve_0_targ_lt_axi_m_wlast(o_pve_0_targ_lt_axi_m_wlast),
        .i_pve_0_targ_lt_axi_m_wready(i_pve_0_targ_lt_axi_m_wready),
        .o_pve_0_targ_lt_axi_m_wstrb(o_pve_0_targ_lt_axi_m_wstrb),
        .o_pve_0_targ_lt_axi_m_wvalid(o_pve_0_targ_lt_axi_m_wvalid),
        .o_pve_0_targ_syscfg_apb_m_paddr(o_pve_0_targ_syscfg_apb_m_paddr),
        .o_pve_0_targ_syscfg_apb_m_penable(o_pve_0_targ_syscfg_apb_m_penable),
        .o_pve_0_targ_syscfg_apb_m_pprot(o_pve_0_targ_syscfg_apb_m_pprot),
        .i_pve_0_targ_syscfg_apb_m_prdata(i_pve_0_targ_syscfg_apb_m_prdata),
        .i_pve_0_targ_syscfg_apb_m_pready(i_pve_0_targ_syscfg_apb_m_pready),
        .o_pve_0_targ_syscfg_apb_m_psel(o_pve_0_targ_syscfg_apb_m_psel),
        .i_pve_0_targ_syscfg_apb_m_pslverr(i_pve_0_targ_syscfg_apb_m_pslverr),
        .o_pve_0_targ_syscfg_apb_m_pstrb(o_pve_0_targ_syscfg_apb_m_pstrb),
        .o_pve_0_targ_syscfg_apb_m_pwdata(o_pve_0_targ_syscfg_apb_m_pwdata),
        .o_pve_0_targ_syscfg_apb_m_pwrite(o_pve_0_targ_syscfg_apb_m_pwrite),
        .i_pve_1_aon_clk(i_pve_1_aon_clk),
        .i_pve_1_aon_rst_n(i_pve_1_aon_rst_n),
        .i_pve_1_clk(i_pve_1_clk),
        .i_pve_1_clken(i_pve_1_clken),
        .i_pve_1_init_ht_axi_s_araddr(i_pve_1_init_ht_axi_s_araddr),
        .i_pve_1_init_ht_axi_s_arburst(i_pve_1_init_ht_axi_s_arburst),
        .i_pve_1_init_ht_axi_s_arcache(i_pve_1_init_ht_axi_s_arcache),
        .i_pve_1_init_ht_axi_s_arid(i_pve_1_init_ht_axi_s_arid),
        .i_pve_1_init_ht_axi_s_arlen(i_pve_1_init_ht_axi_s_arlen),
        .i_pve_1_init_ht_axi_s_arlock(i_pve_1_init_ht_axi_s_arlock),
        .i_pve_1_init_ht_axi_s_arprot(i_pve_1_init_ht_axi_s_arprot),
        .o_pve_1_init_ht_axi_s_arready(o_pve_1_init_ht_axi_s_arready),
        .i_pve_1_init_ht_axi_s_arsize(i_pve_1_init_ht_axi_s_arsize),
        .i_pve_1_init_ht_axi_s_arvalid(i_pve_1_init_ht_axi_s_arvalid),
        .o_pve_1_init_ht_axi_s_rdata(o_pve_1_init_ht_axi_s_rdata),
        .o_pve_1_init_ht_axi_s_rid(o_pve_1_init_ht_axi_s_rid),
        .o_pve_1_init_ht_axi_s_rlast(o_pve_1_init_ht_axi_s_rlast),
        .i_pve_1_init_ht_axi_s_rready(i_pve_1_init_ht_axi_s_rready),
        .o_pve_1_init_ht_axi_s_rresp(o_pve_1_init_ht_axi_s_rresp),
        .o_pve_1_init_ht_axi_s_rvalid(o_pve_1_init_ht_axi_s_rvalid),
        .i_pve_1_init_ht_axi_s_awaddr(i_pve_1_init_ht_axi_s_awaddr),
        .i_pve_1_init_ht_axi_s_awburst(i_pve_1_init_ht_axi_s_awburst),
        .i_pve_1_init_ht_axi_s_awcache(i_pve_1_init_ht_axi_s_awcache),
        .i_pve_1_init_ht_axi_s_awid(i_pve_1_init_ht_axi_s_awid),
        .i_pve_1_init_ht_axi_s_awlen(i_pve_1_init_ht_axi_s_awlen),
        .i_pve_1_init_ht_axi_s_awlock(i_pve_1_init_ht_axi_s_awlock),
        .i_pve_1_init_ht_axi_s_awprot(i_pve_1_init_ht_axi_s_awprot),
        .o_pve_1_init_ht_axi_s_awready(o_pve_1_init_ht_axi_s_awready),
        .i_pve_1_init_ht_axi_s_awsize(i_pve_1_init_ht_axi_s_awsize),
        .i_pve_1_init_ht_axi_s_awvalid(i_pve_1_init_ht_axi_s_awvalid),
        .o_pve_1_init_ht_axi_s_bid(o_pve_1_init_ht_axi_s_bid),
        .i_pve_1_init_ht_axi_s_bready(i_pve_1_init_ht_axi_s_bready),
        .o_pve_1_init_ht_axi_s_bresp(o_pve_1_init_ht_axi_s_bresp),
        .o_pve_1_init_ht_axi_s_bvalid(o_pve_1_init_ht_axi_s_bvalid),
        .i_pve_1_init_ht_axi_s_wdata(i_pve_1_init_ht_axi_s_wdata),
        .i_pve_1_init_ht_axi_s_wlast(i_pve_1_init_ht_axi_s_wlast),
        .o_pve_1_init_ht_axi_s_wready(o_pve_1_init_ht_axi_s_wready),
        .i_pve_1_init_ht_axi_s_wstrb(i_pve_1_init_ht_axi_s_wstrb),
        .i_pve_1_init_ht_axi_s_wvalid(i_pve_1_init_ht_axi_s_wvalid),
        .i_pve_1_init_lt_axi_s_araddr(i_pve_1_init_lt_axi_s_araddr),
        .i_pve_1_init_lt_axi_s_arburst(i_pve_1_init_lt_axi_s_arburst),
        .i_pve_1_init_lt_axi_s_arcache(i_pve_1_init_lt_axi_s_arcache),
        .i_pve_1_init_lt_axi_s_arid(i_pve_1_init_lt_axi_s_arid),
        .i_pve_1_init_lt_axi_s_arlen(i_pve_1_init_lt_axi_s_arlen),
        .i_pve_1_init_lt_axi_s_arlock(i_pve_1_init_lt_axi_s_arlock),
        .i_pve_1_init_lt_axi_s_arprot(i_pve_1_init_lt_axi_s_arprot),
        .i_pve_1_init_lt_axi_s_arqos(i_pve_1_init_lt_axi_s_arqos),
        .o_pve_1_init_lt_axi_s_arready(o_pve_1_init_lt_axi_s_arready),
        .i_pve_1_init_lt_axi_s_arsize(i_pve_1_init_lt_axi_s_arsize),
        .i_pve_1_init_lt_axi_s_arvalid(i_pve_1_init_lt_axi_s_arvalid),
        .o_pve_1_init_lt_axi_s_rdata(o_pve_1_init_lt_axi_s_rdata),
        .o_pve_1_init_lt_axi_s_rid(o_pve_1_init_lt_axi_s_rid),
        .o_pve_1_init_lt_axi_s_rlast(o_pve_1_init_lt_axi_s_rlast),
        .i_pve_1_init_lt_axi_s_rready(i_pve_1_init_lt_axi_s_rready),
        .o_pve_1_init_lt_axi_s_rresp(o_pve_1_init_lt_axi_s_rresp),
        .o_pve_1_init_lt_axi_s_rvalid(o_pve_1_init_lt_axi_s_rvalid),
        .i_pve_1_init_lt_axi_s_awaddr(i_pve_1_init_lt_axi_s_awaddr),
        .i_pve_1_init_lt_axi_s_awburst(i_pve_1_init_lt_axi_s_awburst),
        .i_pve_1_init_lt_axi_s_awcache(i_pve_1_init_lt_axi_s_awcache),
        .i_pve_1_init_lt_axi_s_awid(i_pve_1_init_lt_axi_s_awid),
        .i_pve_1_init_lt_axi_s_awlen(i_pve_1_init_lt_axi_s_awlen),
        .i_pve_1_init_lt_axi_s_awlock(i_pve_1_init_lt_axi_s_awlock),
        .i_pve_1_init_lt_axi_s_awprot(i_pve_1_init_lt_axi_s_awprot),
        .i_pve_1_init_lt_axi_s_awqos(i_pve_1_init_lt_axi_s_awqos),
        .o_pve_1_init_lt_axi_s_awready(o_pve_1_init_lt_axi_s_awready),
        .i_pve_1_init_lt_axi_s_awsize(i_pve_1_init_lt_axi_s_awsize),
        .i_pve_1_init_lt_axi_s_awvalid(i_pve_1_init_lt_axi_s_awvalid),
        .o_pve_1_init_lt_axi_s_bid(o_pve_1_init_lt_axi_s_bid),
        .i_pve_1_init_lt_axi_s_bready(i_pve_1_init_lt_axi_s_bready),
        .o_pve_1_init_lt_axi_s_bresp(o_pve_1_init_lt_axi_s_bresp),
        .o_pve_1_init_lt_axi_s_bvalid(o_pve_1_init_lt_axi_s_bvalid),
        .i_pve_1_init_lt_axi_s_wdata(i_pve_1_init_lt_axi_s_wdata),
        .i_pve_1_init_lt_axi_s_wlast(i_pve_1_init_lt_axi_s_wlast),
        .o_pve_1_init_lt_axi_s_wready(o_pve_1_init_lt_axi_s_wready),
        .i_pve_1_init_lt_axi_s_wstrb(i_pve_1_init_lt_axi_s_wstrb),
        .i_pve_1_init_lt_axi_s_wvalid(i_pve_1_init_lt_axi_s_wvalid),
        .o_pve_1_pwr_idle_val(o_pve_1_pwr_idle_val),
        .o_pve_1_pwr_idle_ack(o_pve_1_pwr_idle_ack),
        .i_pve_1_pwr_idle_req(i_pve_1_pwr_idle_req),
        .i_pve_1_rst_n(i_pve_1_rst_n),
        .o_pve_1_targ_lt_axi_m_araddr(o_pve_1_targ_lt_axi_m_araddr),
        .o_pve_1_targ_lt_axi_m_arburst(o_pve_1_targ_lt_axi_m_arburst),
        .o_pve_1_targ_lt_axi_m_arcache(o_pve_1_targ_lt_axi_m_arcache),
        .o_pve_1_targ_lt_axi_m_arid(o_pve_1_targ_lt_axi_m_arid),
        .o_pve_1_targ_lt_axi_m_arlen(o_pve_1_targ_lt_axi_m_arlen),
        .o_pve_1_targ_lt_axi_m_arlock(o_pve_1_targ_lt_axi_m_arlock),
        .o_pve_1_targ_lt_axi_m_arprot(o_pve_1_targ_lt_axi_m_arprot),
        .o_pve_1_targ_lt_axi_m_arqos(o_pve_1_targ_lt_axi_m_arqos),
        .i_pve_1_targ_lt_axi_m_arready(i_pve_1_targ_lt_axi_m_arready),
        .o_pve_1_targ_lt_axi_m_arsize(o_pve_1_targ_lt_axi_m_arsize),
        .o_pve_1_targ_lt_axi_m_arvalid(o_pve_1_targ_lt_axi_m_arvalid),
        .o_pve_1_targ_lt_axi_m_awaddr(o_pve_1_targ_lt_axi_m_awaddr),
        .o_pve_1_targ_lt_axi_m_awburst(o_pve_1_targ_lt_axi_m_awburst),
        .o_pve_1_targ_lt_axi_m_awcache(o_pve_1_targ_lt_axi_m_awcache),
        .o_pve_1_targ_lt_axi_m_awid(o_pve_1_targ_lt_axi_m_awid),
        .o_pve_1_targ_lt_axi_m_awlen(o_pve_1_targ_lt_axi_m_awlen),
        .o_pve_1_targ_lt_axi_m_awlock(o_pve_1_targ_lt_axi_m_awlock),
        .o_pve_1_targ_lt_axi_m_awprot(o_pve_1_targ_lt_axi_m_awprot),
        .o_pve_1_targ_lt_axi_m_awqos(o_pve_1_targ_lt_axi_m_awqos),
        .i_pve_1_targ_lt_axi_m_awready(i_pve_1_targ_lt_axi_m_awready),
        .o_pve_1_targ_lt_axi_m_awsize(o_pve_1_targ_lt_axi_m_awsize),
        .o_pve_1_targ_lt_axi_m_awvalid(o_pve_1_targ_lt_axi_m_awvalid),
        .i_pve_1_targ_lt_axi_m_bid(i_pve_1_targ_lt_axi_m_bid),
        .o_pve_1_targ_lt_axi_m_bready(o_pve_1_targ_lt_axi_m_bready),
        .i_pve_1_targ_lt_axi_m_bresp(i_pve_1_targ_lt_axi_m_bresp),
        .i_pve_1_targ_lt_axi_m_bvalid(i_pve_1_targ_lt_axi_m_bvalid),
        .i_pve_1_targ_lt_axi_m_rdata(i_pve_1_targ_lt_axi_m_rdata),
        .i_pve_1_targ_lt_axi_m_rid(i_pve_1_targ_lt_axi_m_rid),
        .i_pve_1_targ_lt_axi_m_rlast(i_pve_1_targ_lt_axi_m_rlast),
        .o_pve_1_targ_lt_axi_m_rready(o_pve_1_targ_lt_axi_m_rready),
        .i_pve_1_targ_lt_axi_m_rresp(i_pve_1_targ_lt_axi_m_rresp),
        .i_pve_1_targ_lt_axi_m_rvalid(i_pve_1_targ_lt_axi_m_rvalid),
        .o_pve_1_targ_lt_axi_m_wdata(o_pve_1_targ_lt_axi_m_wdata),
        .o_pve_1_targ_lt_axi_m_wlast(o_pve_1_targ_lt_axi_m_wlast),
        .i_pve_1_targ_lt_axi_m_wready(i_pve_1_targ_lt_axi_m_wready),
        .o_pve_1_targ_lt_axi_m_wstrb(o_pve_1_targ_lt_axi_m_wstrb),
        .o_pve_1_targ_lt_axi_m_wvalid(o_pve_1_targ_lt_axi_m_wvalid),
        .o_pve_1_targ_syscfg_apb_m_paddr(o_pve_1_targ_syscfg_apb_m_paddr),
        .o_pve_1_targ_syscfg_apb_m_penable(o_pve_1_targ_syscfg_apb_m_penable),
        .o_pve_1_targ_syscfg_apb_m_pprot(o_pve_1_targ_syscfg_apb_m_pprot),
        .i_pve_1_targ_syscfg_apb_m_prdata(i_pve_1_targ_syscfg_apb_m_prdata),
        .i_pve_1_targ_syscfg_apb_m_pready(i_pve_1_targ_syscfg_apb_m_pready),
        .o_pve_1_targ_syscfg_apb_m_psel(o_pve_1_targ_syscfg_apb_m_psel),
        .i_pve_1_targ_syscfg_apb_m_pslverr(i_pve_1_targ_syscfg_apb_m_pslverr),
        .o_pve_1_targ_syscfg_apb_m_pstrb(o_pve_1_targ_syscfg_apb_m_pstrb),
        .o_pve_1_targ_syscfg_apb_m_pwdata(o_pve_1_targ_syscfg_apb_m_pwdata),
        .o_pve_1_targ_syscfg_apb_m_pwrite(o_pve_1_targ_syscfg_apb_m_pwrite),
        .i_soc_mgmt_aon_clk(i_soc_mgmt_aon_clk),
        .i_soc_mgmt_aon_rst_n(i_soc_mgmt_aon_rst_n),
        .i_soc_mgmt_clk(i_soc_mgmt_clk),
        .i_soc_mgmt_clken(i_soc_mgmt_clken),
        .i_soc_mgmt_init_lt_axi_s_araddr(i_soc_mgmt_init_lt_axi_s_araddr),
        .i_soc_mgmt_init_lt_axi_s_arburst(i_soc_mgmt_init_lt_axi_s_arburst),
        .i_soc_mgmt_init_lt_axi_s_arcache(i_soc_mgmt_init_lt_axi_s_arcache),
        .i_soc_mgmt_init_lt_axi_s_arid(i_soc_mgmt_init_lt_axi_s_arid),
        .i_soc_mgmt_init_lt_axi_s_arlen(i_soc_mgmt_init_lt_axi_s_arlen),
        .i_soc_mgmt_init_lt_axi_s_arlock(i_soc_mgmt_init_lt_axi_s_arlock),
        .i_soc_mgmt_init_lt_axi_s_arprot(i_soc_mgmt_init_lt_axi_s_arprot),
        .i_soc_mgmt_init_lt_axi_s_arqos(i_soc_mgmt_init_lt_axi_s_arqos),
        .o_soc_mgmt_init_lt_axi_s_arready(o_soc_mgmt_init_lt_axi_s_arready),
        .i_soc_mgmt_init_lt_axi_s_arsize(i_soc_mgmt_init_lt_axi_s_arsize),
        .i_soc_mgmt_init_lt_axi_s_arvalid(i_soc_mgmt_init_lt_axi_s_arvalid),
        .i_soc_mgmt_init_lt_axi_s_awaddr(i_soc_mgmt_init_lt_axi_s_awaddr),
        .i_soc_mgmt_init_lt_axi_s_awburst(i_soc_mgmt_init_lt_axi_s_awburst),
        .i_soc_mgmt_init_lt_axi_s_awcache(i_soc_mgmt_init_lt_axi_s_awcache),
        .i_soc_mgmt_init_lt_axi_s_awid(i_soc_mgmt_init_lt_axi_s_awid),
        .i_soc_mgmt_init_lt_axi_s_awlen(i_soc_mgmt_init_lt_axi_s_awlen),
        .i_soc_mgmt_init_lt_axi_s_awlock(i_soc_mgmt_init_lt_axi_s_awlock),
        .i_soc_mgmt_init_lt_axi_s_awprot(i_soc_mgmt_init_lt_axi_s_awprot),
        .i_soc_mgmt_init_lt_axi_s_awqos(i_soc_mgmt_init_lt_axi_s_awqos),
        .o_soc_mgmt_init_lt_axi_s_awready(o_soc_mgmt_init_lt_axi_s_awready),
        .i_soc_mgmt_init_lt_axi_s_awsize(i_soc_mgmt_init_lt_axi_s_awsize),
        .i_soc_mgmt_init_lt_axi_s_awvalid(i_soc_mgmt_init_lt_axi_s_awvalid),
        .o_soc_mgmt_init_lt_axi_s_bid(o_soc_mgmt_init_lt_axi_s_bid),
        .i_soc_mgmt_init_lt_axi_s_bready(i_soc_mgmt_init_lt_axi_s_bready),
        .o_soc_mgmt_init_lt_axi_s_bresp(o_soc_mgmt_init_lt_axi_s_bresp),
        .o_soc_mgmt_init_lt_axi_s_bvalid(o_soc_mgmt_init_lt_axi_s_bvalid),
        .o_soc_mgmt_init_lt_axi_s_rdata(o_soc_mgmt_init_lt_axi_s_rdata),
        .o_soc_mgmt_init_lt_axi_s_rid(o_soc_mgmt_init_lt_axi_s_rid),
        .o_soc_mgmt_init_lt_axi_s_rlast(o_soc_mgmt_init_lt_axi_s_rlast),
        .i_soc_mgmt_init_lt_axi_s_rready(i_soc_mgmt_init_lt_axi_s_rready),
        .o_soc_mgmt_init_lt_axi_s_rresp(o_soc_mgmt_init_lt_axi_s_rresp),
        .o_soc_mgmt_init_lt_axi_s_rvalid(o_soc_mgmt_init_lt_axi_s_rvalid),
        .i_soc_mgmt_init_lt_axi_s_wdata(i_soc_mgmt_init_lt_axi_s_wdata),
        .i_soc_mgmt_init_lt_axi_s_wlast(i_soc_mgmt_init_lt_axi_s_wlast),
        .o_soc_mgmt_init_lt_axi_s_wready(o_soc_mgmt_init_lt_axi_s_wready),
        .i_soc_mgmt_init_lt_axi_s_wstrb(i_soc_mgmt_init_lt_axi_s_wstrb),
        .i_soc_mgmt_init_lt_axi_s_wvalid(i_soc_mgmt_init_lt_axi_s_wvalid),
        .o_soc_mgmt_pwr_idle_val(o_soc_mgmt_pwr_idle_val),
        .o_soc_mgmt_pwr_idle_ack(o_soc_mgmt_pwr_idle_ack),
        .i_soc_mgmt_pwr_idle_req(i_soc_mgmt_pwr_idle_req),
        .i_soc_mgmt_rst_n(i_soc_mgmt_rst_n),
        .o_soc_mgmt_targ_lt_axi_m_araddr(o_soc_mgmt_targ_lt_axi_m_araddr),
        .o_soc_mgmt_targ_lt_axi_m_arburst(o_soc_mgmt_targ_lt_axi_m_arburst),
        .o_soc_mgmt_targ_lt_axi_m_arcache(o_soc_mgmt_targ_lt_axi_m_arcache),
        .o_soc_mgmt_targ_lt_axi_m_arid(o_soc_mgmt_targ_lt_axi_m_arid),
        .o_soc_mgmt_targ_lt_axi_m_arlen(o_soc_mgmt_targ_lt_axi_m_arlen),
        .o_soc_mgmt_targ_lt_axi_m_arlock(o_soc_mgmt_targ_lt_axi_m_arlock),
        .o_soc_mgmt_targ_lt_axi_m_arprot(o_soc_mgmt_targ_lt_axi_m_arprot),
        .o_soc_mgmt_targ_lt_axi_m_arqos(o_soc_mgmt_targ_lt_axi_m_arqos),
        .i_soc_mgmt_targ_lt_axi_m_arready(i_soc_mgmt_targ_lt_axi_m_arready),
        .o_soc_mgmt_targ_lt_axi_m_arsize(o_soc_mgmt_targ_lt_axi_m_arsize),
        .o_soc_mgmt_targ_lt_axi_m_arvalid(o_soc_mgmt_targ_lt_axi_m_arvalid),
        .o_soc_mgmt_targ_lt_axi_m_awaddr(o_soc_mgmt_targ_lt_axi_m_awaddr),
        .o_soc_mgmt_targ_lt_axi_m_awburst(o_soc_mgmt_targ_lt_axi_m_awburst),
        .o_soc_mgmt_targ_lt_axi_m_awcache(o_soc_mgmt_targ_lt_axi_m_awcache),
        .o_soc_mgmt_targ_lt_axi_m_awid(o_soc_mgmt_targ_lt_axi_m_awid),
        .o_soc_mgmt_targ_lt_axi_m_awlen(o_soc_mgmt_targ_lt_axi_m_awlen),
        .o_soc_mgmt_targ_lt_axi_m_awlock(o_soc_mgmt_targ_lt_axi_m_awlock),
        .o_soc_mgmt_targ_lt_axi_m_awprot(o_soc_mgmt_targ_lt_axi_m_awprot),
        .o_soc_mgmt_targ_lt_axi_m_awqos(o_soc_mgmt_targ_lt_axi_m_awqos),
        .i_soc_mgmt_targ_lt_axi_m_awready(i_soc_mgmt_targ_lt_axi_m_awready),
        .o_soc_mgmt_targ_lt_axi_m_awsize(o_soc_mgmt_targ_lt_axi_m_awsize),
        .o_soc_mgmt_targ_lt_axi_m_awvalid(o_soc_mgmt_targ_lt_axi_m_awvalid),
        .i_soc_mgmt_targ_lt_axi_m_bid(i_soc_mgmt_targ_lt_axi_m_bid),
        .o_soc_mgmt_targ_lt_axi_m_bready(o_soc_mgmt_targ_lt_axi_m_bready),
        .i_soc_mgmt_targ_lt_axi_m_bresp(i_soc_mgmt_targ_lt_axi_m_bresp),
        .i_soc_mgmt_targ_lt_axi_m_bvalid(i_soc_mgmt_targ_lt_axi_m_bvalid),
        .i_soc_mgmt_targ_lt_axi_m_rdata(i_soc_mgmt_targ_lt_axi_m_rdata),
        .i_soc_mgmt_targ_lt_axi_m_rid(i_soc_mgmt_targ_lt_axi_m_rid),
        .i_soc_mgmt_targ_lt_axi_m_rlast(i_soc_mgmt_targ_lt_axi_m_rlast),
        .o_soc_mgmt_targ_lt_axi_m_rready(o_soc_mgmt_targ_lt_axi_m_rready),
        .i_soc_mgmt_targ_lt_axi_m_rresp(i_soc_mgmt_targ_lt_axi_m_rresp),
        .i_soc_mgmt_targ_lt_axi_m_rvalid(i_soc_mgmt_targ_lt_axi_m_rvalid),
        .o_soc_mgmt_targ_lt_axi_m_wdata(o_soc_mgmt_targ_lt_axi_m_wdata),
        .o_soc_mgmt_targ_lt_axi_m_wlast(o_soc_mgmt_targ_lt_axi_m_wlast),
        .i_soc_mgmt_targ_lt_axi_m_wready(i_soc_mgmt_targ_lt_axi_m_wready),
        .o_soc_mgmt_targ_lt_axi_m_wstrb(o_soc_mgmt_targ_lt_axi_m_wstrb),
        .o_soc_mgmt_targ_lt_axi_m_wvalid(o_soc_mgmt_targ_lt_axi_m_wvalid),
        .o_soc_mgmt_targ_syscfg_apb_m_paddr(o_soc_mgmt_targ_syscfg_apb_m_paddr),
        .o_soc_mgmt_targ_syscfg_apb_m_penable(o_soc_mgmt_targ_syscfg_apb_m_penable),
        .o_soc_mgmt_targ_syscfg_apb_m_pprot(o_soc_mgmt_targ_syscfg_apb_m_pprot),
        .i_soc_mgmt_targ_syscfg_apb_m_prdata(i_soc_mgmt_targ_syscfg_apb_m_prdata),
        .i_soc_mgmt_targ_syscfg_apb_m_pready(i_soc_mgmt_targ_syscfg_apb_m_pready),
        .o_soc_mgmt_targ_syscfg_apb_m_psel(o_soc_mgmt_targ_syscfg_apb_m_psel),
        .i_soc_mgmt_targ_syscfg_apb_m_pslverr(i_soc_mgmt_targ_syscfg_apb_m_pslverr),
        .o_soc_mgmt_targ_syscfg_apb_m_pstrb(o_soc_mgmt_targ_syscfg_apb_m_pstrb),
        .o_soc_mgmt_targ_syscfg_apb_m_pwdata(o_soc_mgmt_targ_syscfg_apb_m_pwdata),
        .o_soc_mgmt_targ_syscfg_apb_m_pwrite(o_soc_mgmt_targ_syscfg_apb_m_pwrite),
        .i_sys_spm_aon_clk(i_sys_spm_aon_clk),
        .i_sys_spm_aon_rst_n(i_sys_spm_aon_rst_n),
        .i_sys_spm_clk(i_sys_spm_clk),
        .i_sys_spm_clken(i_sys_spm_clken),
        .o_sys_spm_pwr_idle_val(o_sys_spm_pwr_idle_val),
        .o_sys_spm_pwr_idle_ack(o_sys_spm_pwr_idle_ack),
        .i_sys_spm_pwr_idle_req(i_sys_spm_pwr_idle_req),
        .i_sys_spm_rst_n(i_sys_spm_rst_n),
        .o_sys_spm_targ_lt_axi_m_araddr(o_sys_spm_targ_lt_axi_m_araddr),
        .o_sys_spm_targ_lt_axi_m_arburst(o_sys_spm_targ_lt_axi_m_arburst),
        .o_sys_spm_targ_lt_axi_m_arcache(o_sys_spm_targ_lt_axi_m_arcache),
        .o_sys_spm_targ_lt_axi_m_arid(o_sys_spm_targ_lt_axi_m_arid),
        .o_sys_spm_targ_lt_axi_m_arlen(o_sys_spm_targ_lt_axi_m_arlen),
        .o_sys_spm_targ_lt_axi_m_arlock(o_sys_spm_targ_lt_axi_m_arlock),
        .o_sys_spm_targ_lt_axi_m_arprot(o_sys_spm_targ_lt_axi_m_arprot),
        .o_sys_spm_targ_lt_axi_m_arqos(o_sys_spm_targ_lt_axi_m_arqos),
        .i_sys_spm_targ_lt_axi_m_arready(i_sys_spm_targ_lt_axi_m_arready),
        .o_sys_spm_targ_lt_axi_m_arsize(o_sys_spm_targ_lt_axi_m_arsize),
        .o_sys_spm_targ_lt_axi_m_arvalid(o_sys_spm_targ_lt_axi_m_arvalid),
        .o_sys_spm_targ_lt_axi_m_awaddr(o_sys_spm_targ_lt_axi_m_awaddr),
        .o_sys_spm_targ_lt_axi_m_awburst(o_sys_spm_targ_lt_axi_m_awburst),
        .o_sys_spm_targ_lt_axi_m_awcache(o_sys_spm_targ_lt_axi_m_awcache),
        .o_sys_spm_targ_lt_axi_m_awid(o_sys_spm_targ_lt_axi_m_awid),
        .o_sys_spm_targ_lt_axi_m_awlen(o_sys_spm_targ_lt_axi_m_awlen),
        .o_sys_spm_targ_lt_axi_m_awlock(o_sys_spm_targ_lt_axi_m_awlock),
        .o_sys_spm_targ_lt_axi_m_awprot(o_sys_spm_targ_lt_axi_m_awprot),
        .o_sys_spm_targ_lt_axi_m_awqos(o_sys_spm_targ_lt_axi_m_awqos),
        .i_sys_spm_targ_lt_axi_m_awready(i_sys_spm_targ_lt_axi_m_awready),
        .o_sys_spm_targ_lt_axi_m_awsize(o_sys_spm_targ_lt_axi_m_awsize),
        .o_sys_spm_targ_lt_axi_m_awvalid(o_sys_spm_targ_lt_axi_m_awvalid),
        .i_sys_spm_targ_lt_axi_m_bid(i_sys_spm_targ_lt_axi_m_bid),
        .o_sys_spm_targ_lt_axi_m_bready(o_sys_spm_targ_lt_axi_m_bready),
        .i_sys_spm_targ_lt_axi_m_bresp(i_sys_spm_targ_lt_axi_m_bresp),
        .i_sys_spm_targ_lt_axi_m_bvalid(i_sys_spm_targ_lt_axi_m_bvalid),
        .i_sys_spm_targ_lt_axi_m_rdata(i_sys_spm_targ_lt_axi_m_rdata),
        .i_sys_spm_targ_lt_axi_m_rid(i_sys_spm_targ_lt_axi_m_rid),
        .i_sys_spm_targ_lt_axi_m_rlast(i_sys_spm_targ_lt_axi_m_rlast),
        .o_sys_spm_targ_lt_axi_m_rready(o_sys_spm_targ_lt_axi_m_rready),
        .i_sys_spm_targ_lt_axi_m_rresp(i_sys_spm_targ_lt_axi_m_rresp),
        .i_sys_spm_targ_lt_axi_m_rvalid(i_sys_spm_targ_lt_axi_m_rvalid),
        .o_sys_spm_targ_lt_axi_m_wdata(o_sys_spm_targ_lt_axi_m_wdata),
        .o_sys_spm_targ_lt_axi_m_wlast(o_sys_spm_targ_lt_axi_m_wlast),
        .i_sys_spm_targ_lt_axi_m_wready(i_sys_spm_targ_lt_axi_m_wready),
        .o_sys_spm_targ_lt_axi_m_wstrb(o_sys_spm_targ_lt_axi_m_wstrb),
        .o_sys_spm_targ_lt_axi_m_wvalid(o_sys_spm_targ_lt_axi_m_wvalid),
        .o_sys_spm_targ_syscfg_apb_m_paddr(o_sys_spm_targ_syscfg_apb_m_paddr),
        .o_sys_spm_targ_syscfg_apb_m_penable(o_sys_spm_targ_syscfg_apb_m_penable),
        .o_sys_spm_targ_syscfg_apb_m_pprot(o_sys_spm_targ_syscfg_apb_m_pprot),
        .i_sys_spm_targ_syscfg_apb_m_prdata(i_sys_spm_targ_syscfg_apb_m_prdata),
        .i_sys_spm_targ_syscfg_apb_m_pready(i_sys_spm_targ_syscfg_apb_m_pready),
        .o_sys_spm_targ_syscfg_apb_m_psel(o_sys_spm_targ_syscfg_apb_m_psel),
        .i_sys_spm_targ_syscfg_apb_m_pslverr(i_sys_spm_targ_syscfg_apb_m_pslverr),
        .o_sys_spm_targ_syscfg_apb_m_pstrb(o_sys_spm_targ_syscfg_apb_m_pstrb),
        .o_sys_spm_targ_syscfg_apb_m_pwdata(o_sys_spm_targ_syscfg_apb_m_pwdata),
        .o_sys_spm_targ_syscfg_apb_m_pwrite(o_sys_spm_targ_syscfg_apb_m_pwrite),

        // Token Network IOs
        // -- NIUs
        .i_apu_init_tok_ocpl_s_maddr(i_apu_init_tok_ocpl_s_maddr),
        .i_apu_init_tok_ocpl_s_mcmd(i_apu_init_tok_ocpl_s_mcmd),
        .i_apu_init_tok_ocpl_s_mdata(i_apu_init_tok_ocpl_s_mdata),
        .o_apu_init_tok_ocpl_s_scmdaccept(o_apu_init_tok_ocpl_s_scmdaccept),
        .o_apu_pwr_tok_idle_val(o_apu_pwr_tok_idle_val),
        .o_apu_pwr_tok_idle_ack(o_apu_pwr_tok_idle_ack),
        .i_apu_pwr_tok_idle_req(i_apu_pwr_tok_idle_req),
        .o_apu_targ_tok_ocpl_m_maddr(o_apu_targ_tok_ocpl_m_maddr),
        .o_apu_targ_tok_ocpl_m_mcmd(o_apu_targ_tok_ocpl_m_mcmd),
        .o_apu_targ_tok_ocpl_m_mdata(o_apu_targ_tok_ocpl_m_mdata),
        .i_apu_targ_tok_ocpl_m_scmdaccept(i_apu_targ_tok_ocpl_m_scmdaccept),

        .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_data),
        .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_head),
        .o_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_rdy),
        .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_tail),
        .i_dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld(dp_lnk_cross_east_to_soc_tok_0_egress_to_lnk_cross_east_to_soc_tok_0_ingress_vld),
        .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_data),
        .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_head),
        .o_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_rdy),
        .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_tail),
        .i_dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld(dp_lnk_cross_east_to_soc_tok_1_egress_to_lnk_cross_east_to_soc_tok_1_ingress_vld),
        .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_data),
        .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_head),
        .i_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_rdy),
        .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_tail),
        .o_dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld(dp_lnk_cross_soc_to_east_tok_0_egress_to_lnk_cross_soc_to_east_tok_0_ingress_vld),
        .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_data),
        .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_head),
        .i_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_rdy),
        .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_tail),
        .o_dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld(dp_lnk_cross_soc_to_east_tok_1_egress_to_lnk_cross_soc_to_east_tok_1_ingress_vld),

        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  ),
        .bisr_clk('0),
        .bisr_reset('0),
        .bisr_shift_en('0),
        .bisr_si('0),
        .bisr_so(  )
    );

    chip_pkg::chip_syscfg_addr_t            center_to_sdma_0_cfg_apb4_paddr;
    chip_pkg::chip_apb_syscfg_data_t        center_to_sdma_0_cfg_apb4_pwdata;
    logic                                   center_to_sdma_0_cfg_apb4_pwrite;
    logic                                   center_to_sdma_0_cfg_apb4_psel;
    logic                                   center_to_sdma_0_cfg_apb4_penable;
    chip_pkg::chip_apb_syscfg_strb_t        center_to_sdma_0_cfg_apb4_pstrb;
    logic [3-1:0]                           center_to_sdma_0_cfg_apb4_pprot;
    logic                                   center_to_sdma_0_cfg_apb4_pready;
    chip_pkg::chip_apb_syscfg_data_t        center_to_sdma_0_cfg_apb4_prdata;
    logic                                   center_to_sdma_0_cfg_apb4_pslverr;
    logic                                   center_to_sdma_0_noc_async_idle_req;
    logic                                   center_to_sdma_0_noc_async_idle_ack;
    logic                                   center_to_sdma_0_noc_async_idle_val;
    logic                                   center_to_sdma_0_noc_tok_async_idle_req;
    logic                                   center_to_sdma_0_noc_tok_async_idle_ack;
    logic                                   center_to_sdma_0_noc_tok_async_idle_val;
    logic                                   center_to_sdma_0_noc_clken;
    logic                                   center_to_sdma_0_noc_rst_n;
    logic                                   center_to_sdma_0_targ_lt_axi_awvalid;
    chip_pkg::chip_axi_addr_t               center_to_sdma_0_targ_lt_axi_awaddr;
    sdma_pkg::sdma_axi_lt_id_t              center_to_sdma_0_targ_lt_axi_awid;
    axi_pkg::axi_len_t                      center_to_sdma_0_targ_lt_axi_awlen;
    axi_pkg::axi_size_t                     center_to_sdma_0_targ_lt_axi_awsize;
    axi_pkg::axi_burst_t                    center_to_sdma_0_targ_lt_axi_awburst;
    logic                                   center_to_sdma_0_targ_lt_axi_awlock;
    axi_pkg::axi_cache_t                    center_to_sdma_0_targ_lt_axi_awcache;
    axi_pkg::axi_prot_t                     center_to_sdma_0_targ_lt_axi_awprot;
    logic                                   center_to_sdma_0_targ_lt_axi_awready;
    logic                                   center_to_sdma_0_targ_lt_axi_wvalid;
    logic                                   center_to_sdma_0_targ_lt_axi_wlast;
    chip_pkg::chip_axi_lt_data_t            center_to_sdma_0_targ_lt_axi_wdata;
    chip_pkg::chip_axi_lt_wstrb_t           center_to_sdma_0_targ_lt_axi_wstrb;
    logic                                   center_to_sdma_0_targ_lt_axi_wready;
    logic                                   center_to_sdma_0_targ_lt_axi_bvalid;
    sdma_pkg::sdma_axi_lt_id_t              center_to_sdma_0_targ_lt_axi_bid;
    axi_pkg::axi_resp_e                     center_to_sdma_0_targ_lt_axi_bresp;
    logic                                   center_to_sdma_0_targ_lt_axi_bready;
    logic                                   center_to_sdma_0_targ_lt_axi_arvalid;
    chip_pkg::chip_axi_addr_t               center_to_sdma_0_targ_lt_axi_araddr;
    sdma_pkg::sdma_axi_lt_id_t              center_to_sdma_0_targ_lt_axi_arid;
    axi_pkg::axi_len_t                      center_to_sdma_0_targ_lt_axi_arlen;
    axi_pkg::axi_size_t                     center_to_sdma_0_targ_lt_axi_arsize;
    axi_pkg::axi_burst_t                    center_to_sdma_0_targ_lt_axi_arburst;
    logic                                   center_to_sdma_0_targ_lt_axi_arlock;
    axi_pkg::axi_cache_t                    center_to_sdma_0_targ_lt_axi_arcache;
    axi_pkg::axi_prot_t                     center_to_sdma_0_targ_lt_axi_arprot;
    logic                                   center_to_sdma_0_targ_lt_axi_arready;
    logic                                   center_to_sdma_0_targ_lt_axi_rvalid;
    logic                                   center_to_sdma_0_targ_lt_axi_rlast;
    sdma_pkg::sdma_axi_lt_id_t              center_to_sdma_0_targ_lt_axi_rid;
    chip_pkg::chip_axi_lt_data_t            center_to_sdma_0_targ_lt_axi_rdata;
    axi_pkg::axi_resp_e                     center_to_sdma_0_targ_lt_axi_rresp;
    logic                                   center_to_sdma_0_targ_lt_axi_rready;
    logic                                   sdma_0_to_center_init_ht_0_axi_awvalid;
    chip_pkg::chip_axi_addr_t               sdma_0_to_center_init_ht_0_axi_awaddr;
    sdma_pkg::sdma_axi_ht_id_t              sdma_0_to_center_init_ht_0_axi_awid;
    axi_pkg::axi_len_t                      sdma_0_to_center_init_ht_0_axi_awlen;
    axi_pkg::axi_size_e                     sdma_0_to_center_init_ht_0_axi_awsize;
    axi_pkg::axi_burst_e                    sdma_0_to_center_init_ht_0_axi_awburst;
    logic                                   sdma_0_to_center_init_ht_0_axi_awlock;
    axi_pkg::axi_cache_e                    sdma_0_to_center_init_ht_0_axi_awcache;
    axi_pkg::axi_prot_t                     sdma_0_to_center_init_ht_0_axi_awprot;
    logic                                   sdma_0_to_center_init_ht_0_axi_awready;
    logic                                   sdma_0_to_center_init_ht_0_axi_wvalid;
    logic                                   sdma_0_to_center_init_ht_0_axi_wlast;
    chip_pkg::chip_axi_ht_data_t            sdma_0_to_center_init_ht_0_axi_wdata;
    chip_pkg::chip_axi_ht_wstrb_t           sdma_0_to_center_init_ht_0_axi_wstrb;
    logic                                   sdma_0_to_center_init_ht_0_axi_wready;
    logic                                   sdma_0_to_center_init_ht_0_axi_bvalid;
    sdma_pkg::sdma_axi_ht_id_t              sdma_0_to_center_init_ht_0_axi_bid;
    axi_pkg::axi_resp_t                     sdma_0_to_center_init_ht_0_axi_bresp;
    logic                                   sdma_0_to_center_init_ht_0_axi_bready;
    logic                                   sdma_0_to_center_init_ht_0_axi_arvalid;
    chip_pkg::chip_axi_addr_t               sdma_0_to_center_init_ht_0_axi_araddr;
    sdma_pkg::sdma_axi_ht_id_t              sdma_0_to_center_init_ht_0_axi_arid;
    axi_pkg::axi_len_t                      sdma_0_to_center_init_ht_0_axi_arlen;
    axi_pkg::axi_size_e                     sdma_0_to_center_init_ht_0_axi_arsize;
    axi_pkg::axi_burst_e                    sdma_0_to_center_init_ht_0_axi_arburst;
    logic                                   sdma_0_to_center_init_ht_0_axi_arlock;
    axi_pkg::axi_cache_e                    sdma_0_to_center_init_ht_0_axi_arcache;
    axi_pkg::axi_prot_t                     sdma_0_to_center_init_ht_0_axi_arprot;
    logic                                   sdma_0_to_center_init_ht_0_axi_arready;
    logic                                   sdma_0_to_center_init_ht_0_axi_rvalid;
    logic                                   sdma_0_to_center_init_ht_0_axi_rlast;
    sdma_pkg::sdma_axi_ht_id_t              sdma_0_to_center_init_ht_0_axi_rid;
    chip_pkg::chip_axi_ht_data_t            sdma_0_to_center_init_ht_0_axi_rdata;
    axi_pkg::axi_resp_t                     sdma_0_to_center_init_ht_0_axi_rresp;
    logic                                   sdma_0_to_center_init_ht_0_axi_rready;
    logic                                   sdma_0_to_center_init_ht_1_axi_awvalid;
    chip_pkg::chip_axi_addr_t               sdma_0_to_center_init_ht_1_axi_awaddr;
    sdma_pkg::sdma_axi_ht_id_t              sdma_0_to_center_init_ht_1_axi_awid;
    axi_pkg::axi_len_t                      sdma_0_to_center_init_ht_1_axi_awlen;
    axi_pkg::axi_size_e                     sdma_0_to_center_init_ht_1_axi_awsize;
    axi_pkg::axi_burst_e                    sdma_0_to_center_init_ht_1_axi_awburst;
    logic                                   sdma_0_to_center_init_ht_1_axi_awlock;
    axi_pkg::axi_cache_e                    sdma_0_to_center_init_ht_1_axi_awcache;
    axi_pkg::axi_prot_t                     sdma_0_to_center_init_ht_1_axi_awprot;
    logic                                   sdma_0_to_center_init_ht_1_axi_awready;
    logic                                   sdma_0_to_center_init_ht_1_axi_wvalid;
    logic                                   sdma_0_to_center_init_ht_1_axi_wlast;
    chip_pkg::chip_axi_ht_data_t            sdma_0_to_center_init_ht_1_axi_wdata;
    chip_pkg::chip_axi_ht_wstrb_t           sdma_0_to_center_init_ht_1_axi_wstrb;
    logic                                   sdma_0_to_center_init_ht_1_axi_wready;
    logic                                   sdma_0_to_center_init_ht_1_axi_bvalid;
    sdma_pkg::sdma_axi_ht_id_t              sdma_0_to_center_init_ht_1_axi_bid;
    axi_pkg::axi_resp_t                     sdma_0_to_center_init_ht_1_axi_bresp;
    logic                                   sdma_0_to_center_init_ht_1_axi_bready;
    logic                                   sdma_0_to_center_init_ht_1_axi_arvalid;
    chip_pkg::chip_axi_addr_t               sdma_0_to_center_init_ht_1_axi_araddr;
    sdma_pkg::sdma_axi_ht_id_t              sdma_0_to_center_init_ht_1_axi_arid;
    axi_pkg::axi_len_t                      sdma_0_to_center_init_ht_1_axi_arlen;
    axi_pkg::axi_size_e                     sdma_0_to_center_init_ht_1_axi_arsize;
    axi_pkg::axi_burst_e                    sdma_0_to_center_init_ht_1_axi_arburst;
    logic                                   sdma_0_to_center_init_ht_1_axi_arlock;
    axi_pkg::axi_cache_e                    sdma_0_to_center_init_ht_1_axi_arcache;
    axi_pkg::axi_prot_t                     sdma_0_to_center_init_ht_1_axi_arprot;
    logic                                   sdma_0_to_center_init_ht_1_axi_arready;
    logic                                   sdma_0_to_center_init_ht_1_axi_rvalid;
    logic                                   sdma_0_to_center_init_ht_1_axi_rlast;
    sdma_pkg::sdma_axi_ht_id_t              sdma_0_to_center_init_ht_1_axi_rid;
    chip_pkg::chip_axi_ht_data_t            sdma_0_to_center_init_ht_1_axi_rdata;
    axi_pkg::axi_resp_t                     sdma_0_to_center_init_ht_1_axi_rresp;
    logic                                   sdma_0_to_center_init_ht_1_axi_rready;
    sdma_pkg::sdma_axi_lt_id_t              sdma_0_to_center_init_lt_awid;
    chip_pkg::chip_axi_addr_t               sdma_0_to_center_init_lt_awaddr;
    axi_pkg::axi_len_t                      sdma_0_to_center_init_lt_awlen;
    axi_pkg::axi_size_t                     sdma_0_to_center_init_lt_awsize;
    axi_pkg::axi_burst_t                    sdma_0_to_center_init_lt_awburst;
    axi_pkg::axi_cache_t                    sdma_0_to_center_init_lt_awcache;
    axi_pkg::axi_qos_t                      sdma_0_to_center_init_lt_awqos;
    logic                                   sdma_0_to_center_init_lt_awlock;
    axi_pkg::axi_prot_t                     sdma_0_to_center_init_lt_awprot;
    logic                                   sdma_0_to_center_init_lt_awvalid;
    logic                                   sdma_0_to_center_init_lt_awready;
    chip_pkg::chip_axi_lt_data_t            sdma_0_to_center_init_lt_wdata;
    chip_pkg::chip_axi_lt_wstrb_t           sdma_0_to_center_init_lt_wstrb;
    logic                                   sdma_0_to_center_init_lt_wlast;
    logic                                   sdma_0_to_center_init_lt_wvalid;
    logic                                   sdma_0_to_center_init_lt_wready;
    sdma_pkg::sdma_axi_lt_id_t              sdma_0_to_center_init_lt_bid;
    axi_pkg::axi_resp_t                     sdma_0_to_center_init_lt_bresp;
    logic                                   sdma_0_to_center_init_lt_bvalid;
    logic                                   sdma_0_to_center_init_lt_bready;
    sdma_pkg::sdma_axi_lt_id_t              sdma_0_to_center_init_lt_arid;
    chip_pkg::chip_axi_addr_t               sdma_0_to_center_init_lt_araddr;
    axi_pkg::axi_len_t                      sdma_0_to_center_init_lt_arlen;
    axi_pkg::axi_size_t                     sdma_0_to_center_init_lt_arsize;
    axi_pkg::axi_burst_t                    sdma_0_to_center_init_lt_arburst;
    axi_pkg::axi_cache_t                    sdma_0_to_center_init_lt_arcache;
    axi_pkg::axi_qos_t                      sdma_0_to_center_init_lt_arqos;
    logic                                   sdma_0_to_center_init_lt_arlock;
    axi_pkg::axi_prot_t                     sdma_0_to_center_init_lt_arprot;
    logic                                   sdma_0_to_center_init_lt_arvalid;
    logic                                   sdma_0_to_center_init_lt_arready;
    sdma_pkg::sdma_axi_lt_id_t              sdma_0_to_center_init_lt_rid;
    chip_pkg::chip_axi_lt_data_t            sdma_0_to_center_init_lt_rdata;
    axi_pkg::axi_resp_t                     sdma_0_to_center_init_lt_rresp;
    logic                                   sdma_0_to_center_init_lt_rlast;
    logic                                   sdma_0_to_center_init_lt_rvalid;
    logic                                   sdma_0_to_center_init_lt_rready;

    chip_pkg::chip_syscfg_addr_t            center_to_sdma_1_cfg_apb4_paddr;
    chip_pkg::chip_apb_syscfg_data_t        center_to_sdma_1_cfg_apb4_pwdata;
    logic                                   center_to_sdma_1_cfg_apb4_pwrite;
    logic                                   center_to_sdma_1_cfg_apb4_psel;
    logic                                   center_to_sdma_1_cfg_apb4_penable;
    chip_pkg::chip_apb_syscfg_strb_t        center_to_sdma_1_cfg_apb4_pstrb;
    logic [3-1:0]                           center_to_sdma_1_cfg_apb4_pprot;
    logic                                   center_to_sdma_1_cfg_apb4_pready;
    chip_pkg::chip_apb_syscfg_data_t        center_to_sdma_1_cfg_apb4_prdata;
    logic                                   center_to_sdma_1_cfg_apb4_pslverr;
    logic                                   center_to_sdma_1_noc_async_idle_req;
    logic                                   center_to_sdma_1_noc_async_idle_ack;
    logic                                   center_to_sdma_1_noc_async_idle_val;
    logic                                   center_to_sdma_1_noc_tok_async_idle_req;
    logic                                   center_to_sdma_1_noc_tok_async_idle_ack;
    logic                                   center_to_sdma_1_noc_tok_async_idle_val;
    logic                                   center_to_sdma_1_noc_clken;
    logic                                   center_to_sdma_1_noc_rst_n;
    logic                                   center_to_sdma_1_targ_lt_axi_awvalid;
    chip_pkg::chip_axi_addr_t               center_to_sdma_1_targ_lt_axi_awaddr;
    sdma_pkg::sdma_axi_lt_id_t              center_to_sdma_1_targ_lt_axi_awid;
    axi_pkg::axi_len_t                      center_to_sdma_1_targ_lt_axi_awlen;
    axi_pkg::axi_size_t                     center_to_sdma_1_targ_lt_axi_awsize;
    axi_pkg::axi_burst_t                    center_to_sdma_1_targ_lt_axi_awburst;
    logic                                   center_to_sdma_1_targ_lt_axi_awlock;
    axi_pkg::axi_cache_t                    center_to_sdma_1_targ_lt_axi_awcache;
    axi_pkg::axi_prot_t                     center_to_sdma_1_targ_lt_axi_awprot;
    logic                                   center_to_sdma_1_targ_lt_axi_awready;
    logic                                   center_to_sdma_1_targ_lt_axi_wvalid;
    logic                                   center_to_sdma_1_targ_lt_axi_wlast;
    chip_pkg::chip_axi_lt_data_t            center_to_sdma_1_targ_lt_axi_wdata;
    chip_pkg::chip_axi_lt_wstrb_t           center_to_sdma_1_targ_lt_axi_wstrb;
    logic                                   center_to_sdma_1_targ_lt_axi_wready;
    logic                                   center_to_sdma_1_targ_lt_axi_bvalid;
    sdma_pkg::sdma_axi_lt_id_t              center_to_sdma_1_targ_lt_axi_bid;
    axi_pkg::axi_resp_e                     center_to_sdma_1_targ_lt_axi_bresp;
    logic                                   center_to_sdma_1_targ_lt_axi_bready;
    logic                                   center_to_sdma_1_targ_lt_axi_arvalid;
    chip_pkg::chip_axi_addr_t               center_to_sdma_1_targ_lt_axi_araddr;
    sdma_pkg::sdma_axi_lt_id_t              center_to_sdma_1_targ_lt_axi_arid;
    axi_pkg::axi_len_t                      center_to_sdma_1_targ_lt_axi_arlen;
    axi_pkg::axi_size_t                     center_to_sdma_1_targ_lt_axi_arsize;
    axi_pkg::axi_burst_t                    center_to_sdma_1_targ_lt_axi_arburst;
    logic                                   center_to_sdma_1_targ_lt_axi_arlock;
    axi_pkg::axi_cache_t                    center_to_sdma_1_targ_lt_axi_arcache;
    axi_pkg::axi_prot_t                     center_to_sdma_1_targ_lt_axi_arprot;
    logic                                   center_to_sdma_1_targ_lt_axi_arready;
    logic                                   center_to_sdma_1_targ_lt_axi_rvalid;
    logic                                   center_to_sdma_1_targ_lt_axi_rlast;
    sdma_pkg::sdma_axi_lt_id_t              center_to_sdma_1_targ_lt_axi_rid;
    chip_pkg::chip_axi_lt_data_t            center_to_sdma_1_targ_lt_axi_rdata;
    axi_pkg::axi_resp_e                     center_to_sdma_1_targ_lt_axi_rresp;
    logic                                   center_to_sdma_1_targ_lt_axi_rready;
    logic                                   sdma_1_to_center_init_ht_0_axi_awvalid;
    chip_pkg::chip_axi_addr_t               sdma_1_to_center_init_ht_0_axi_awaddr;
    sdma_pkg::sdma_axi_ht_id_t              sdma_1_to_center_init_ht_0_axi_awid;
    axi_pkg::axi_len_t                      sdma_1_to_center_init_ht_0_axi_awlen;
    axi_pkg::axi_size_e                     sdma_1_to_center_init_ht_0_axi_awsize;
    axi_pkg::axi_burst_e                    sdma_1_to_center_init_ht_0_axi_awburst;
    logic                                   sdma_1_to_center_init_ht_0_axi_awlock;
    axi_pkg::axi_cache_e                    sdma_1_to_center_init_ht_0_axi_awcache;
    axi_pkg::axi_prot_t                     sdma_1_to_center_init_ht_0_axi_awprot;
    logic                                   sdma_1_to_center_init_ht_0_axi_awready;
    logic                                   sdma_1_to_center_init_ht_0_axi_wvalid;
    logic                                   sdma_1_to_center_init_ht_0_axi_wlast;
    chip_pkg::chip_axi_ht_data_t            sdma_1_to_center_init_ht_0_axi_wdata;
    chip_pkg::chip_axi_ht_wstrb_t           sdma_1_to_center_init_ht_0_axi_wstrb;
    logic                                   sdma_1_to_center_init_ht_0_axi_wready;
    logic                                   sdma_1_to_center_init_ht_0_axi_bvalid;
    sdma_pkg::sdma_axi_ht_id_t              sdma_1_to_center_init_ht_0_axi_bid;
    axi_pkg::axi_resp_t                     sdma_1_to_center_init_ht_0_axi_bresp;
    logic                                   sdma_1_to_center_init_ht_0_axi_bready;
    logic                                   sdma_1_to_center_init_ht_0_axi_arvalid;
    chip_pkg::chip_axi_addr_t               sdma_1_to_center_init_ht_0_axi_araddr;
    sdma_pkg::sdma_axi_ht_id_t              sdma_1_to_center_init_ht_0_axi_arid;
    axi_pkg::axi_len_t                      sdma_1_to_center_init_ht_0_axi_arlen;
    axi_pkg::axi_size_e                     sdma_1_to_center_init_ht_0_axi_arsize;
    axi_pkg::axi_burst_e                    sdma_1_to_center_init_ht_0_axi_arburst;
    logic                                   sdma_1_to_center_init_ht_0_axi_arlock;
    axi_pkg::axi_cache_e                    sdma_1_to_center_init_ht_0_axi_arcache;
    axi_pkg::axi_prot_t                     sdma_1_to_center_init_ht_0_axi_arprot;
    logic                                   sdma_1_to_center_init_ht_0_axi_arready;
    logic                                   sdma_1_to_center_init_ht_0_axi_rvalid;
    logic                                   sdma_1_to_center_init_ht_0_axi_rlast;
    sdma_pkg::sdma_axi_ht_id_t              sdma_1_to_center_init_ht_0_axi_rid;
    chip_pkg::chip_axi_ht_data_t            sdma_1_to_center_init_ht_0_axi_rdata;
    axi_pkg::axi_resp_t                     sdma_1_to_center_init_ht_0_axi_rresp;
    logic                                   sdma_1_to_center_init_ht_0_axi_rready;
    logic                                   sdma_1_to_center_init_ht_1_axi_awvalid;
    chip_pkg::chip_axi_addr_t               sdma_1_to_center_init_ht_1_axi_awaddr;
    sdma_pkg::sdma_axi_ht_id_t              sdma_1_to_center_init_ht_1_axi_awid;
    axi_pkg::axi_len_t                      sdma_1_to_center_init_ht_1_axi_awlen;
    axi_pkg::axi_size_e                     sdma_1_to_center_init_ht_1_axi_awsize;
    axi_pkg::axi_burst_e                    sdma_1_to_center_init_ht_1_axi_awburst;
    logic                                   sdma_1_to_center_init_ht_1_axi_awlock;
    axi_pkg::axi_cache_e                    sdma_1_to_center_init_ht_1_axi_awcache;
    axi_pkg::axi_prot_t                     sdma_1_to_center_init_ht_1_axi_awprot;
    logic                                   sdma_1_to_center_init_ht_1_axi_awready;
    logic                                   sdma_1_to_center_init_ht_1_axi_wvalid;
    logic                                   sdma_1_to_center_init_ht_1_axi_wlast;
    chip_pkg::chip_axi_ht_data_t            sdma_1_to_center_init_ht_1_axi_wdata;
    chip_pkg::chip_axi_ht_wstrb_t           sdma_1_to_center_init_ht_1_axi_wstrb;
    logic                                   sdma_1_to_center_init_ht_1_axi_wready;
    logic                                   sdma_1_to_center_init_ht_1_axi_bvalid;
    sdma_pkg::sdma_axi_ht_id_t              sdma_1_to_center_init_ht_1_axi_bid;
    axi_pkg::axi_resp_t                     sdma_1_to_center_init_ht_1_axi_bresp;
    logic                                   sdma_1_to_center_init_ht_1_axi_bready;
    logic                                   sdma_1_to_center_init_ht_1_axi_arvalid;
    chip_pkg::chip_axi_addr_t               sdma_1_to_center_init_ht_1_axi_araddr;
    sdma_pkg::sdma_axi_ht_id_t              sdma_1_to_center_init_ht_1_axi_arid;
    axi_pkg::axi_len_t                      sdma_1_to_center_init_ht_1_axi_arlen;
    axi_pkg::axi_size_e                     sdma_1_to_center_init_ht_1_axi_arsize;
    axi_pkg::axi_burst_e                    sdma_1_to_center_init_ht_1_axi_arburst;
    logic                                   sdma_1_to_center_init_ht_1_axi_arlock;
    axi_pkg::axi_cache_e                    sdma_1_to_center_init_ht_1_axi_arcache;
    axi_pkg::axi_prot_t                     sdma_1_to_center_init_ht_1_axi_arprot;
    logic                                   sdma_1_to_center_init_ht_1_axi_arready;
    logic                                   sdma_1_to_center_init_ht_1_axi_rvalid;
    logic                                   sdma_1_to_center_init_ht_1_axi_rlast;
    sdma_pkg::sdma_axi_ht_id_t              sdma_1_to_center_init_ht_1_axi_rid;
    chip_pkg::chip_axi_ht_data_t            sdma_1_to_center_init_ht_1_axi_rdata;
    axi_pkg::axi_resp_t                     sdma_1_to_center_init_ht_1_axi_rresp;
    logic                                   sdma_1_to_center_init_ht_1_axi_rready;
    sdma_pkg::sdma_axi_lt_id_t              sdma_1_to_center_init_lt_awid;
    chip_pkg::chip_axi_addr_t               sdma_1_to_center_init_lt_awaddr;
    axi_pkg::axi_len_t                      sdma_1_to_center_init_lt_awlen;
    axi_pkg::axi_size_t                     sdma_1_to_center_init_lt_awsize;
    axi_pkg::axi_burst_t                    sdma_1_to_center_init_lt_awburst;
    axi_pkg::axi_cache_t                    sdma_1_to_center_init_lt_awcache;
    axi_pkg::axi_qos_t                      sdma_1_to_center_init_lt_awqos;
    logic                                   sdma_1_to_center_init_lt_awlock;
    axi_pkg::axi_prot_t                     sdma_1_to_center_init_lt_awprot;
    logic                                   sdma_1_to_center_init_lt_awvalid;
    logic                                   sdma_1_to_center_init_lt_awready;
    chip_pkg::chip_axi_lt_data_t            sdma_1_to_center_init_lt_wdata;
    chip_pkg::chip_axi_lt_wstrb_t           sdma_1_to_center_init_lt_wstrb;
    logic                                   sdma_1_to_center_init_lt_wlast;
    logic                                   sdma_1_to_center_init_lt_wvalid;
    logic                                   sdma_1_to_center_init_lt_wready;
    sdma_pkg::sdma_axi_lt_id_t              sdma_1_to_center_init_lt_bid;
    axi_pkg::axi_resp_t                     sdma_1_to_center_init_lt_bresp;
    logic                                   sdma_1_to_center_init_lt_bvalid;
    logic                                   sdma_1_to_center_init_lt_bready;
    sdma_pkg::sdma_axi_lt_id_t              sdma_1_to_center_init_lt_arid;
    chip_pkg::chip_axi_addr_t               sdma_1_to_center_init_lt_araddr;
    axi_pkg::axi_len_t                      sdma_1_to_center_init_lt_arlen;
    axi_pkg::axi_size_t                     sdma_1_to_center_init_lt_arsize;
    axi_pkg::axi_burst_t                    sdma_1_to_center_init_lt_arburst;
    axi_pkg::axi_cache_t                    sdma_1_to_center_init_lt_arcache;
    axi_pkg::axi_qos_t                      sdma_1_to_center_init_lt_arqos;
    logic                                   sdma_1_to_center_init_lt_arlock;
    axi_pkg::axi_prot_t                     sdma_1_to_center_init_lt_arprot;
    logic                                   sdma_1_to_center_init_lt_arvalid;
    logic                                   sdma_1_to_center_init_lt_arready;
    sdma_pkg::sdma_axi_lt_id_t              sdma_1_to_center_init_lt_rid;
    chip_pkg::chip_axi_lt_data_t            sdma_1_to_center_init_lt_rdata;
    axi_pkg::axi_resp_t                     sdma_1_to_center_init_lt_rresp;
    logic                                   sdma_1_to_center_init_lt_rlast;
    logic                                   sdma_1_to_center_init_lt_rvalid;
    logic                                   sdma_1_to_center_init_lt_rready;

    // SDMA 0
    logic                             sdma_0_init_tok_ocpl_mcmd;
    logic                             sdma_0_init_tok_ocpl_scmdaccept;
    chip_pkg::chip_ocpl_token_addr_t  sdma_0_init_tok_ocpl_maddr;
    chip_pkg::chip_ocpl_token_data_t  sdma_0_init_tok_ocpl_mdata;
    chip_pkg::chip_ocpl_token_addr_t  sdma_0_targ_tok_ocpl_maddr;
    logic                             sdma_0_targ_tok_ocpl_mcmd;
    logic                             sdma_0_targ_tok_ocpl_scmdaccept;
    chip_pkg::chip_ocpl_token_data_t  sdma_0_targ_tok_ocpl_mdata;

    sdma_p u_sdma_0_p(
        .i_clk             (i_sdma_0_clk),
        .i_ref_clk         (i_ref_clk),
        .i_ao_rst_n        (i_sdma_0_ao_rst_n),
        .i_global_rst_n    (i_sdma_0_global_rst_n),
        .o_int             (o_sdma_0_int),
        .i_sdma_nr         (1'b0),
        .i_inter_core_sync (i_sdma_inter_core_sync),

        // Token Network
        .o_tok_prod_ocpl_m_maddr      (sdma_0_init_tok_ocpl_maddr),
        .o_tok_prod_ocpl_m_mcmd       (sdma_0_init_tok_ocpl_mcmd),
        .i_tok_prod_ocpl_m_scmdaccept (sdma_0_init_tok_ocpl_scmdaccept),
        .o_tok_prod_ocpl_m_mdata      (sdma_0_init_tok_ocpl_mdata),
        .i_tok_cons_ocpl_s_maddr      (sdma_0_targ_tok_ocpl_maddr),
        .i_tok_cons_ocpl_s_mcmd       (sdma_0_targ_tok_ocpl_mcmd),
        .o_tok_cons_ocpl_s_scmdaccept (sdma_0_targ_tok_ocpl_scmdaccept),
        .i_tok_cons_ocpl_s_mdata      (sdma_0_targ_tok_ocpl_mdata),
        .o_noc_tok_async_idle_req     (center_to_sdma_0_noc_tok_async_idle_req),
        .i_noc_tok_async_idle_ack     (center_to_sdma_0_noc_tok_async_idle_ack),
        .i_noc_tok_async_idle_val     (center_to_sdma_0_noc_tok_async_idle_val),

        .i_cfg_apb4_s_paddr         (center_to_sdma_0_cfg_apb4_paddr),
        .i_cfg_apb4_s_pwdata        (center_to_sdma_0_cfg_apb4_pwdata),
        .i_cfg_apb4_s_pwrite        (center_to_sdma_0_cfg_apb4_pwrite),
        .i_cfg_apb4_s_psel          (center_to_sdma_0_cfg_apb4_psel),
        .i_cfg_apb4_s_penable       (center_to_sdma_0_cfg_apb4_penable),
        .i_cfg_apb4_s_pstrb         (center_to_sdma_0_cfg_apb4_pstrb),
        .i_cfg_apb4_s_pprot         (center_to_sdma_0_cfg_apb4_pprot),
        .o_cfg_apb4_s_pready        (center_to_sdma_0_cfg_apb4_pready),
        .o_cfg_apb4_s_prdata        (center_to_sdma_0_cfg_apb4_prdata),
        .o_cfg_apb4_s_pslverr       (center_to_sdma_0_cfg_apb4_pslverr),
        .o_noc_async_idle_req       (center_to_sdma_0_noc_async_idle_req),
        .i_noc_async_idle_ack       (center_to_sdma_0_noc_async_idle_ack),
        .i_noc_async_idle_val       (center_to_sdma_0_noc_async_idle_val),
        .o_noc_clken                (center_to_sdma_0_noc_clken),
        .o_noc_rst_n                (center_to_sdma_0_noc_rst_n),
        .i_clock_throttle           (i_sdma_0_clock_throttle),
        .i_axi_s_awvalid            (center_to_sdma_0_targ_lt_axi_awvalid),
        .i_axi_s_awaddr             (center_to_sdma_0_targ_lt_axi_awaddr),
        .i_axi_s_awid               (center_to_sdma_0_targ_lt_axi_awid),
        .i_axi_s_awlen              (center_to_sdma_0_targ_lt_axi_awlen),
        .i_axi_s_awsize             (axi_pkg::axi_size_e'(center_to_sdma_0_targ_lt_axi_awsize)),
        .i_axi_s_awburst            (axi_pkg::axi_burst_e'(center_to_sdma_0_targ_lt_axi_awburst)),
        .i_axi_s_awlock             (center_to_sdma_0_targ_lt_axi_awlock),
        .i_axi_s_awcache            (axi_pkg::axi_cache_e'(center_to_sdma_0_targ_lt_axi_awcache)),
        .i_axi_s_awprot             (center_to_sdma_0_targ_lt_axi_awprot),
        .o_axi_s_awready            (center_to_sdma_0_targ_lt_axi_awready),
        .i_axi_s_wvalid             (center_to_sdma_0_targ_lt_axi_wvalid),
        .i_axi_s_wlast              (center_to_sdma_0_targ_lt_axi_wlast),
        .i_axi_s_wdata              (center_to_sdma_0_targ_lt_axi_wdata),
        .i_axi_s_wstrb              (center_to_sdma_0_targ_lt_axi_wstrb),
        .o_axi_s_wready             (center_to_sdma_0_targ_lt_axi_wready),
        .o_axi_s_bvalid             (center_to_sdma_0_targ_lt_axi_bvalid),
        .o_axi_s_bid                (center_to_sdma_0_targ_lt_axi_bid),
        .o_axi_s_bresp              (center_to_sdma_0_targ_lt_axi_bresp),
        .i_axi_s_bready             (center_to_sdma_0_targ_lt_axi_bready),
        .i_axi_s_arvalid            (center_to_sdma_0_targ_lt_axi_arvalid),
        .i_axi_s_araddr             (center_to_sdma_0_targ_lt_axi_araddr),
        .i_axi_s_arid               (center_to_sdma_0_targ_lt_axi_arid),
        .i_axi_s_arlen              (center_to_sdma_0_targ_lt_axi_arlen),
        .i_axi_s_arsize             (axi_pkg::axi_size_e'(center_to_sdma_0_targ_lt_axi_arsize)),
        .i_axi_s_arburst            (axi_pkg::axi_burst_e'(center_to_sdma_0_targ_lt_axi_arburst)),
        .i_axi_s_arlock             (center_to_sdma_0_targ_lt_axi_arlock),
        .i_axi_s_arcache            (axi_pkg::axi_cache_e'(center_to_sdma_0_targ_lt_axi_arcache)),
        .i_axi_s_arprot             (center_to_sdma_0_targ_lt_axi_arprot),
        .o_axi_s_arready            (center_to_sdma_0_targ_lt_axi_arready),
        .o_axi_s_rvalid             (center_to_sdma_0_targ_lt_axi_rvalid),
        .o_axi_s_rlast              (center_to_sdma_0_targ_lt_axi_rlast),
        .o_axi_s_rid                (center_to_sdma_0_targ_lt_axi_rid),
        .o_axi_s_rdata              (center_to_sdma_0_targ_lt_axi_rdata),
        .o_axi_s_rresp              (center_to_sdma_0_targ_lt_axi_rresp),
        .i_axi_s_rready             (center_to_sdma_0_targ_lt_axi_rready),
        .o_axi_m0_awvalid           (sdma_0_to_center_init_ht_0_axi_awvalid),
        .o_axi_m0_awaddr            (sdma_0_to_center_init_ht_0_axi_awaddr),
        .o_axi_m0_awid              (sdma_0_to_center_init_ht_0_axi_awid),
        .o_axi_m0_awlen             (sdma_0_to_center_init_ht_0_axi_awlen),
        .o_axi_m0_awsize            (sdma_0_to_center_init_ht_0_axi_awsize),
        .o_axi_m0_awburst           (sdma_0_to_center_init_ht_0_axi_awburst),
        .o_axi_m0_awlock            (sdma_0_to_center_init_ht_0_axi_awlock),
        .o_axi_m0_awcache           (sdma_0_to_center_init_ht_0_axi_awcache),
        .o_axi_m0_awprot            (sdma_0_to_center_init_ht_0_axi_awprot),
        .i_axi_m0_awready           (sdma_0_to_center_init_ht_0_axi_awready),
        .o_axi_m0_wvalid            (sdma_0_to_center_init_ht_0_axi_wvalid),
        .o_axi_m0_wlast             (sdma_0_to_center_init_ht_0_axi_wlast),
        .o_axi_m0_wdata             (sdma_0_to_center_init_ht_0_axi_wdata),
        .o_axi_m0_wstrb             (sdma_0_to_center_init_ht_0_axi_wstrb),
        .i_axi_m0_wready            (sdma_0_to_center_init_ht_0_axi_wready),
        .i_axi_m0_bvalid            (sdma_0_to_center_init_ht_0_axi_bvalid),
        .i_axi_m0_bid               (sdma_0_to_center_init_ht_0_axi_bid),
        .i_axi_m0_bresp             (axi_pkg::axi_resp_e'(sdma_0_to_center_init_ht_0_axi_bresp)),
        .o_axi_m0_bready            (sdma_0_to_center_init_ht_0_axi_bready),
        .o_axi_m0_arvalid           (sdma_0_to_center_init_ht_0_axi_arvalid),
        .o_axi_m0_araddr            (sdma_0_to_center_init_ht_0_axi_araddr),
        .o_axi_m0_arid              (sdma_0_to_center_init_ht_0_axi_arid),
        .o_axi_m0_arlen             (sdma_0_to_center_init_ht_0_axi_arlen),
        .o_axi_m0_arsize            (sdma_0_to_center_init_ht_0_axi_arsize),
        .o_axi_m0_arburst           (sdma_0_to_center_init_ht_0_axi_arburst),
        .o_axi_m0_arlock            (sdma_0_to_center_init_ht_0_axi_arlock),
        .o_axi_m0_arcache           (sdma_0_to_center_init_ht_0_axi_arcache),
        .o_axi_m0_arprot            (sdma_0_to_center_init_ht_0_axi_arprot),
        .i_axi_m0_arready           (sdma_0_to_center_init_ht_0_axi_arready),
        .i_axi_m0_rvalid            (sdma_0_to_center_init_ht_0_axi_rvalid),
        .i_axi_m0_rlast             (sdma_0_to_center_init_ht_0_axi_rlast),
        .i_axi_m0_rid               (sdma_0_to_center_init_ht_0_axi_rid),
        .i_axi_m0_rdata             (sdma_0_to_center_init_ht_0_axi_rdata),
        .i_axi_m0_rresp             (axi_pkg::axi_resp_e'(sdma_0_to_center_init_ht_0_axi_rresp)),
        .o_axi_m0_rready            (sdma_0_to_center_init_ht_0_axi_rready),
        .o_axi_m1_awvalid           (sdma_0_to_center_init_ht_1_axi_awvalid),
        .o_axi_m1_awaddr            (sdma_0_to_center_init_ht_1_axi_awaddr),
        .o_axi_m1_awid              (sdma_0_to_center_init_ht_1_axi_awid),
        .o_axi_m1_awlen             (sdma_0_to_center_init_ht_1_axi_awlen),
        .o_axi_m1_awsize            (sdma_0_to_center_init_ht_1_axi_awsize),
        .o_axi_m1_awburst           (sdma_0_to_center_init_ht_1_axi_awburst),
        .o_axi_m1_awlock            (sdma_0_to_center_init_ht_1_axi_awlock),
        .o_axi_m1_awcache           (sdma_0_to_center_init_ht_1_axi_awcache),
        .o_axi_m1_awprot            (sdma_0_to_center_init_ht_1_axi_awprot),
        .i_axi_m1_awready           (sdma_0_to_center_init_ht_1_axi_awready),
        .o_axi_m1_wvalid            (sdma_0_to_center_init_ht_1_axi_wvalid),
        .o_axi_m1_wlast             (sdma_0_to_center_init_ht_1_axi_wlast),
        .o_axi_m1_wdata             (sdma_0_to_center_init_ht_1_axi_wdata),
        .o_axi_m1_wstrb             (sdma_0_to_center_init_ht_1_axi_wstrb),
        .i_axi_m1_wready            (sdma_0_to_center_init_ht_1_axi_wready),
        .i_axi_m1_bvalid            (sdma_0_to_center_init_ht_1_axi_bvalid),
        .i_axi_m1_bid               (sdma_0_to_center_init_ht_1_axi_bid),
        .i_axi_m1_bresp             (axi_pkg::axi_resp_e'(sdma_0_to_center_init_ht_1_axi_bresp)),
        .o_axi_m1_bready            (sdma_0_to_center_init_ht_1_axi_bready),
        .o_axi_m1_arvalid           (sdma_0_to_center_init_ht_1_axi_arvalid),
        .o_axi_m1_araddr            (sdma_0_to_center_init_ht_1_axi_araddr),
        .o_axi_m1_arid              (sdma_0_to_center_init_ht_1_axi_arid),
        .o_axi_m1_arlen             (sdma_0_to_center_init_ht_1_axi_arlen),
        .o_axi_m1_arsize            (sdma_0_to_center_init_ht_1_axi_arsize),
        .o_axi_m1_arburst           (sdma_0_to_center_init_ht_1_axi_arburst),
        .o_axi_m1_arlock            (sdma_0_to_center_init_ht_1_axi_arlock),
        .o_axi_m1_arcache           (sdma_0_to_center_init_ht_1_axi_arcache),
        .o_axi_m1_arprot            (sdma_0_to_center_init_ht_1_axi_arprot),
        .i_axi_m1_arready           (sdma_0_to_center_init_ht_1_axi_arready),
        .i_axi_m1_rvalid            (sdma_0_to_center_init_ht_1_axi_rvalid),
        .i_axi_m1_rlast             (sdma_0_to_center_init_ht_1_axi_rlast),
        .i_axi_m1_rid               (sdma_0_to_center_init_ht_1_axi_rid),
        .i_axi_m1_rdata             (sdma_0_to_center_init_ht_1_axi_rdata),
        .i_axi_m1_rresp             (axi_pkg::axi_resp_e'(sdma_0_to_center_init_ht_1_axi_rresp)),
        .o_axi_m1_rready            (sdma_0_to_center_init_ht_1_axi_rready),
        .o_axi_trc_m_awid           (sdma_0_to_center_init_lt_awid),
        .o_axi_trc_m_awaddr         (sdma_0_to_center_init_lt_awaddr),
        .o_axi_trc_m_awlen          (sdma_0_to_center_init_lt_awlen),
        .o_axi_trc_m_awsize         (sdma_0_to_center_init_lt_awsize),
        .o_axi_trc_m_awburst        (sdma_0_to_center_init_lt_awburst),
        .o_axi_trc_m_awcache        (sdma_0_to_center_init_lt_awcache),
        .o_axi_trc_m_awlock         (sdma_0_to_center_init_lt_awlock),
        .o_axi_trc_m_awprot         (sdma_0_to_center_init_lt_awprot),
        .o_axi_trc_m_awqos          (sdma_0_to_center_init_lt_awqos),
        .o_axi_trc_m_awvalid        (sdma_0_to_center_init_lt_awvalid),
        .i_axi_trc_m_awready        (sdma_0_to_center_init_lt_awready),
        .o_axi_trc_m_wdata          (sdma_0_to_center_init_lt_wdata),
        .o_axi_trc_m_wstrb          (sdma_0_to_center_init_lt_wstrb),
        .o_axi_trc_m_wlast          (sdma_0_to_center_init_lt_wlast),
        .o_axi_trc_m_wvalid         (sdma_0_to_center_init_lt_wvalid),
        .i_axi_trc_m_wready         (sdma_0_to_center_init_lt_wready),
        .i_axi_trc_m_bid            (sdma_0_to_center_init_lt_bid),
        .i_axi_trc_m_bresp          (sdma_0_to_center_init_lt_bresp),
        .i_axi_trc_m_bvalid         (sdma_0_to_center_init_lt_bvalid),
        .o_axi_trc_m_bready         (sdma_0_to_center_init_lt_bready),
        .o_axi_trc_m_arid           (sdma_0_to_center_init_lt_arid),
        .o_axi_trc_m_araddr         (sdma_0_to_center_init_lt_araddr),
        .o_axi_trc_m_arlen          (sdma_0_to_center_init_lt_arlen),
        .o_axi_trc_m_arsize         (sdma_0_to_center_init_lt_arsize),
        .o_axi_trc_m_arburst        (sdma_0_to_center_init_lt_arburst),
        .o_axi_trc_m_arcache        (sdma_0_to_center_init_lt_arcache),
        .o_axi_trc_m_arlock         (sdma_0_to_center_init_lt_arlock),
        .o_axi_trc_m_arprot         (sdma_0_to_center_init_lt_arprot),
        .o_axi_trc_m_arqos          (sdma_0_to_center_init_lt_arqos),
        .o_axi_trc_m_arvalid        (sdma_0_to_center_init_lt_arvalid),
        .i_axi_trc_m_arready        (sdma_0_to_center_init_lt_arready),
        .i_axi_trc_m_rid            (sdma_0_to_center_init_lt_rid),
        .i_axi_trc_m_rdata          (sdma_0_to_center_init_lt_rdata),
        .i_axi_trc_m_rresp          (sdma_0_to_center_init_lt_rresp),
        .i_axi_trc_m_rlast          (sdma_0_to_center_init_lt_rlast),
        .i_axi_trc_m_rvalid         (sdma_0_to_center_init_lt_rvalid),
        .o_axi_trc_m_rready         (sdma_0_to_center_init_lt_rready),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  ),
        .bisr_clk('0),
        .bisr_reset('0),
        .bisr_shift_en('0),
        .bisr_si('0),
        .bisr_so(  )

    );


    // SDMA 1
    logic                             sdma_1_init_tok_ocpl_mcmd;
    logic                             sdma_1_init_tok_ocpl_scmdaccept;
    chip_pkg::chip_ocpl_token_addr_t  sdma_1_init_tok_ocpl_maddr;
    chip_pkg::chip_ocpl_token_data_t  sdma_1_init_tok_ocpl_mdata;
    chip_pkg::chip_ocpl_token_addr_t  sdma_1_targ_tok_ocpl_maddr;
    logic                             sdma_1_targ_tok_ocpl_mcmd;
    logic                             sdma_1_targ_tok_ocpl_scmdaccept;
    chip_pkg::chip_ocpl_token_data_t  sdma_1_targ_tok_ocpl_mdata;
    sdma_p u_sdma_1_p(
        .i_clk                      (i_sdma_1_clk),
        .i_ref_clk                  (i_ref_clk),
        .i_ao_rst_n                 (i_sdma_1_ao_rst_n),
        .i_global_rst_n             (i_sdma_1_global_rst_n),
        .o_int                      (o_sdma_1_int),
        .i_sdma_nr                  (1'b1),
        .i_inter_core_sync          (i_sdma_inter_core_sync),

        // Token Network
        .o_tok_prod_ocpl_m_maddr      (sdma_1_init_tok_ocpl_maddr),
        .o_tok_prod_ocpl_m_mcmd       (sdma_1_init_tok_ocpl_mcmd),
        .i_tok_prod_ocpl_m_scmdaccept (sdma_1_init_tok_ocpl_scmdaccept),
        .o_tok_prod_ocpl_m_mdata      (sdma_1_init_tok_ocpl_mdata),
        .i_tok_cons_ocpl_s_maddr      (sdma_1_targ_tok_ocpl_maddr),
        .i_tok_cons_ocpl_s_mcmd       (sdma_1_targ_tok_ocpl_mcmd),
        .o_tok_cons_ocpl_s_scmdaccept (sdma_1_targ_tok_ocpl_scmdaccept),
        .i_tok_cons_ocpl_s_mdata      (sdma_1_targ_tok_ocpl_mdata),
        .o_noc_tok_async_idle_req     (center_to_sdma_1_noc_tok_async_idle_req),
        .i_noc_tok_async_idle_ack     (center_to_sdma_1_noc_tok_async_idle_ack),
        .i_noc_tok_async_idle_val     (center_to_sdma_1_noc_tok_async_idle_val),

        .i_cfg_apb4_s_paddr         (center_to_sdma_1_cfg_apb4_paddr),
        .i_cfg_apb4_s_pwdata        (center_to_sdma_1_cfg_apb4_pwdata),
        .i_cfg_apb4_s_pwrite        (center_to_sdma_1_cfg_apb4_pwrite),
        .i_cfg_apb4_s_psel          (center_to_sdma_1_cfg_apb4_psel),
        .i_cfg_apb4_s_penable       (center_to_sdma_1_cfg_apb4_penable),
        .i_cfg_apb4_s_pstrb         (center_to_sdma_1_cfg_apb4_pstrb),
        .i_cfg_apb4_s_pprot         (center_to_sdma_1_cfg_apb4_pprot),
        .o_cfg_apb4_s_pready        (center_to_sdma_1_cfg_apb4_pready),
        .o_cfg_apb4_s_prdata        (center_to_sdma_1_cfg_apb4_prdata),
        .o_cfg_apb4_s_pslverr       (center_to_sdma_1_cfg_apb4_pslverr),
        .o_noc_async_idle_req       (center_to_sdma_1_noc_async_idle_req),
        .i_noc_async_idle_ack       (center_to_sdma_1_noc_async_idle_ack),
        .i_noc_async_idle_val       (center_to_sdma_1_noc_async_idle_val),
        .o_noc_clken                (center_to_sdma_1_noc_clken),
        .o_noc_rst_n                (center_to_sdma_1_noc_rst_n),
        .i_clock_throttle           (i_sdma_1_clock_throttle),
        .i_axi_s_awvalid            (center_to_sdma_1_targ_lt_axi_awvalid),
        .i_axi_s_awaddr             (center_to_sdma_1_targ_lt_axi_awaddr),
        .i_axi_s_awid               (center_to_sdma_1_targ_lt_axi_awid),
        .i_axi_s_awlen              (center_to_sdma_1_targ_lt_axi_awlen),
        .i_axi_s_awsize             (axi_pkg::axi_size_e'(center_to_sdma_1_targ_lt_axi_awsize)),
        .i_axi_s_awburst            (axi_pkg::axi_burst_e'(center_to_sdma_1_targ_lt_axi_awburst)),
        .i_axi_s_awlock             (center_to_sdma_1_targ_lt_axi_awlock),
        .i_axi_s_awcache            (axi_pkg::axi_cache_e'(center_to_sdma_1_targ_lt_axi_awcache)),
        .i_axi_s_awprot             (center_to_sdma_1_targ_lt_axi_awprot),
        .o_axi_s_awready            (center_to_sdma_1_targ_lt_axi_awready),
        .i_axi_s_wvalid             (center_to_sdma_1_targ_lt_axi_wvalid),
        .i_axi_s_wlast              (center_to_sdma_1_targ_lt_axi_wlast),
        .i_axi_s_wdata              (center_to_sdma_1_targ_lt_axi_wdata),
        .i_axi_s_wstrb              (center_to_sdma_1_targ_lt_axi_wstrb),
        .o_axi_s_wready             (center_to_sdma_1_targ_lt_axi_wready),
        .o_axi_s_bvalid             (center_to_sdma_1_targ_lt_axi_bvalid),
        .o_axi_s_bid                (center_to_sdma_1_targ_lt_axi_bid),
        .o_axi_s_bresp              (center_to_sdma_1_targ_lt_axi_bresp),
        .i_axi_s_bready             (center_to_sdma_1_targ_lt_axi_bready),
        .i_axi_s_arvalid            (center_to_sdma_1_targ_lt_axi_arvalid),
        .i_axi_s_araddr             (center_to_sdma_1_targ_lt_axi_araddr),
        .i_axi_s_arid               (center_to_sdma_1_targ_lt_axi_arid),
        .i_axi_s_arlen              (center_to_sdma_1_targ_lt_axi_arlen),
        .i_axi_s_arsize             (axi_pkg::axi_size_e'(center_to_sdma_1_targ_lt_axi_arsize)),
        .i_axi_s_arburst            (axi_pkg::axi_burst_e'(center_to_sdma_1_targ_lt_axi_arburst)),
        .i_axi_s_arlock             (center_to_sdma_1_targ_lt_axi_arlock),
        .i_axi_s_arcache            (axi_pkg::axi_cache_e'(center_to_sdma_1_targ_lt_axi_arcache)),
        .i_axi_s_arprot             (center_to_sdma_1_targ_lt_axi_arprot),
        .o_axi_s_arready            (center_to_sdma_1_targ_lt_axi_arready),
        .o_axi_s_rvalid             (center_to_sdma_1_targ_lt_axi_rvalid),
        .o_axi_s_rlast              (center_to_sdma_1_targ_lt_axi_rlast),
        .o_axi_s_rid                (center_to_sdma_1_targ_lt_axi_rid),
        .o_axi_s_rdata              (center_to_sdma_1_targ_lt_axi_rdata),
        .o_axi_s_rresp              (center_to_sdma_1_targ_lt_axi_rresp),
        .i_axi_s_rready             (center_to_sdma_1_targ_lt_axi_rready),
        .o_axi_m0_awvalid           (sdma_1_to_center_init_ht_0_axi_awvalid),
        .o_axi_m0_awaddr            (sdma_1_to_center_init_ht_0_axi_awaddr),
        .o_axi_m0_awid              (sdma_1_to_center_init_ht_0_axi_awid),
        .o_axi_m0_awlen             (sdma_1_to_center_init_ht_0_axi_awlen),
        .o_axi_m0_awsize            (sdma_1_to_center_init_ht_0_axi_awsize),
        .o_axi_m0_awburst           (sdma_1_to_center_init_ht_0_axi_awburst),
        .o_axi_m0_awlock            (sdma_1_to_center_init_ht_0_axi_awlock),
        .o_axi_m0_awcache           (sdma_1_to_center_init_ht_0_axi_awcache),
        .o_axi_m0_awprot            (sdma_1_to_center_init_ht_0_axi_awprot),
        .i_axi_m0_awready           (sdma_1_to_center_init_ht_0_axi_awready),
        .o_axi_m0_wvalid            (sdma_1_to_center_init_ht_0_axi_wvalid),
        .o_axi_m0_wlast             (sdma_1_to_center_init_ht_0_axi_wlast),
        .o_axi_m0_wdata             (sdma_1_to_center_init_ht_0_axi_wdata),
        .o_axi_m0_wstrb             (sdma_1_to_center_init_ht_0_axi_wstrb),
        .i_axi_m0_wready            (sdma_1_to_center_init_ht_0_axi_wready),
        .i_axi_m0_bvalid            (sdma_1_to_center_init_ht_0_axi_bvalid),
        .i_axi_m0_bid               (sdma_1_to_center_init_ht_0_axi_bid),
        .i_axi_m0_bresp             (axi_pkg::axi_resp_e'(sdma_1_to_center_init_ht_0_axi_bresp)),
        .o_axi_m0_bready            (sdma_1_to_center_init_ht_0_axi_bready),
        .o_axi_m0_arvalid           (sdma_1_to_center_init_ht_0_axi_arvalid),
        .o_axi_m0_araddr            (sdma_1_to_center_init_ht_0_axi_araddr),
        .o_axi_m0_arid              (sdma_1_to_center_init_ht_0_axi_arid),
        .o_axi_m0_arlen             (sdma_1_to_center_init_ht_0_axi_arlen),
        .o_axi_m0_arsize            (sdma_1_to_center_init_ht_0_axi_arsize),
        .o_axi_m0_arburst           (sdma_1_to_center_init_ht_0_axi_arburst),
        .o_axi_m0_arlock            (sdma_1_to_center_init_ht_0_axi_arlock),
        .o_axi_m0_arcache           (sdma_1_to_center_init_ht_0_axi_arcache),
        .o_axi_m0_arprot            (sdma_1_to_center_init_ht_0_axi_arprot),
        .i_axi_m0_arready           (sdma_1_to_center_init_ht_0_axi_arready),
        .i_axi_m0_rvalid            (sdma_1_to_center_init_ht_0_axi_rvalid),
        .i_axi_m0_rlast             (sdma_1_to_center_init_ht_0_axi_rlast),
        .i_axi_m0_rid               (sdma_1_to_center_init_ht_0_axi_rid),
        .i_axi_m0_rdata             (sdma_1_to_center_init_ht_0_axi_rdata),
        .i_axi_m0_rresp             (axi_pkg::axi_resp_e'(sdma_1_to_center_init_ht_0_axi_rresp)),
        .o_axi_m0_rready            (sdma_1_to_center_init_ht_0_axi_rready),
        .o_axi_m1_awvalid           (sdma_1_to_center_init_ht_1_axi_awvalid),
        .o_axi_m1_awaddr            (sdma_1_to_center_init_ht_1_axi_awaddr),
        .o_axi_m1_awid              (sdma_1_to_center_init_ht_1_axi_awid),
        .o_axi_m1_awlen             (sdma_1_to_center_init_ht_1_axi_awlen),
        .o_axi_m1_awsize            (sdma_1_to_center_init_ht_1_axi_awsize),
        .o_axi_m1_awburst           (sdma_1_to_center_init_ht_1_axi_awburst),
        .o_axi_m1_awlock            (sdma_1_to_center_init_ht_1_axi_awlock),
        .o_axi_m1_awcache           (sdma_1_to_center_init_ht_1_axi_awcache),
        .o_axi_m1_awprot            (sdma_1_to_center_init_ht_1_axi_awprot),
        .i_axi_m1_awready           (sdma_1_to_center_init_ht_1_axi_awready),
        .o_axi_m1_wvalid            (sdma_1_to_center_init_ht_1_axi_wvalid),
        .o_axi_m1_wlast             (sdma_1_to_center_init_ht_1_axi_wlast),
        .o_axi_m1_wdata             (sdma_1_to_center_init_ht_1_axi_wdata),
        .o_axi_m1_wstrb             (sdma_1_to_center_init_ht_1_axi_wstrb),
        .i_axi_m1_wready            (sdma_1_to_center_init_ht_1_axi_wready),
        .i_axi_m1_bvalid            (sdma_1_to_center_init_ht_1_axi_bvalid),
        .i_axi_m1_bid               (sdma_1_to_center_init_ht_1_axi_bid),
        .i_axi_m1_bresp             (axi_pkg::axi_resp_e'(sdma_1_to_center_init_ht_1_axi_bresp)),
        .o_axi_m1_bready            (sdma_1_to_center_init_ht_1_axi_bready),
        .o_axi_m1_arvalid           (sdma_1_to_center_init_ht_1_axi_arvalid),
        .o_axi_m1_araddr            (sdma_1_to_center_init_ht_1_axi_araddr),
        .o_axi_m1_arid              (sdma_1_to_center_init_ht_1_axi_arid),
        .o_axi_m1_arlen             (sdma_1_to_center_init_ht_1_axi_arlen),
        .o_axi_m1_arsize            (sdma_1_to_center_init_ht_1_axi_arsize),
        .o_axi_m1_arburst           (sdma_1_to_center_init_ht_1_axi_arburst),
        .o_axi_m1_arlock            (sdma_1_to_center_init_ht_1_axi_arlock),
        .o_axi_m1_arcache           (sdma_1_to_center_init_ht_1_axi_arcache),
        .o_axi_m1_arprot            (sdma_1_to_center_init_ht_1_axi_arprot),
        .i_axi_m1_arready           (sdma_1_to_center_init_ht_1_axi_arready),
        .i_axi_m1_rvalid            (sdma_1_to_center_init_ht_1_axi_rvalid),
        .i_axi_m1_rlast             (sdma_1_to_center_init_ht_1_axi_rlast),
        .i_axi_m1_rid               (sdma_1_to_center_init_ht_1_axi_rid),
        .i_axi_m1_rdata             (sdma_1_to_center_init_ht_1_axi_rdata),
        .i_axi_m1_rresp             (axi_pkg::axi_resp_e'(sdma_1_to_center_init_ht_1_axi_rresp)),
        .o_axi_m1_rready            (sdma_1_to_center_init_ht_1_axi_rready),
        .o_axi_trc_m_awid           (sdma_1_to_center_init_lt_awid),
        .o_axi_trc_m_awaddr         (sdma_1_to_center_init_lt_awaddr),
        .o_axi_trc_m_awlen          (sdma_1_to_center_init_lt_awlen),
        .o_axi_trc_m_awsize         (sdma_1_to_center_init_lt_awsize),
        .o_axi_trc_m_awburst        (sdma_1_to_center_init_lt_awburst),
        .o_axi_trc_m_awcache        (sdma_1_to_center_init_lt_awcache),
        .o_axi_trc_m_awlock         (sdma_1_to_center_init_lt_awlock),
        .o_axi_trc_m_awprot         (sdma_1_to_center_init_lt_awprot),
        .o_axi_trc_m_awqos          (sdma_1_to_center_init_lt_awqos),
        .o_axi_trc_m_awvalid        (sdma_1_to_center_init_lt_awvalid),
        .i_axi_trc_m_awready        (sdma_1_to_center_init_lt_awready),
        .o_axi_trc_m_wdata          (sdma_1_to_center_init_lt_wdata),
        .o_axi_trc_m_wstrb          (sdma_1_to_center_init_lt_wstrb),
        .o_axi_trc_m_wlast          (sdma_1_to_center_init_lt_wlast),
        .o_axi_trc_m_wvalid         (sdma_1_to_center_init_lt_wvalid),
        .i_axi_trc_m_wready         (sdma_1_to_center_init_lt_wready),
        .i_axi_trc_m_bid            (sdma_1_to_center_init_lt_bid),
        .i_axi_trc_m_bresp          (sdma_1_to_center_init_lt_bresp),
        .i_axi_trc_m_bvalid         (sdma_1_to_center_init_lt_bvalid),
        .o_axi_trc_m_bready         (sdma_1_to_center_init_lt_bready),
        .o_axi_trc_m_arid           (sdma_1_to_center_init_lt_arid),
        .o_axi_trc_m_araddr         (sdma_1_to_center_init_lt_araddr),
        .o_axi_trc_m_arlen          (sdma_1_to_center_init_lt_arlen),
        .o_axi_trc_m_arsize         (sdma_1_to_center_init_lt_arsize),
        .o_axi_trc_m_arburst        (sdma_1_to_center_init_lt_arburst),
        .o_axi_trc_m_arcache        (sdma_1_to_center_init_lt_arcache),
        .o_axi_trc_m_arlock         (sdma_1_to_center_init_lt_arlock),
        .o_axi_trc_m_arprot         (sdma_1_to_center_init_lt_arprot),
        .o_axi_trc_m_arqos          (sdma_1_to_center_init_lt_arqos),
        .o_axi_trc_m_arvalid        (sdma_1_to_center_init_lt_arvalid),
        .i_axi_trc_m_arready        (sdma_1_to_center_init_lt_arready),
        .i_axi_trc_m_rid            (sdma_1_to_center_init_lt_rid),
        .i_axi_trc_m_rdata          (sdma_1_to_center_init_lt_rdata),
        .i_axi_trc_m_rresp          (sdma_1_to_center_init_lt_rresp),
        .i_axi_trc_m_rlast          (sdma_1_to_center_init_lt_rlast),
        .i_axi_trc_m_rvalid         (sdma_1_to_center_init_lt_rvalid),
        .o_axi_trc_m_rready         (sdma_1_to_center_init_lt_rready),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  ),
        .bisr_clk('0),
        .bisr_reset('0),
        .bisr_shift_en('0),
        .bisr_si('0),
        .bisr_so(  )

    );

    // Instance of noc_v_center_p
    noc_v_center_p v_center_p (
        .i_sdma_0_aon_clk                       (i_ref_clk),
        .i_sdma_0_aon_rst_n                     (i_sdma_0_ao_rst_n),
        .i_sdma_0_clk                           (i_sdma_0_clk),
        .i_sdma_0_clken                         (center_to_sdma_0_noc_clken),
        .i_sdma_0_init_ht_0_axi_s_araddr        (sdma_0_to_center_init_ht_0_axi_araddr),
        .i_sdma_0_init_ht_0_axi_s_arburst       (sdma_0_to_center_init_ht_0_axi_arburst),
        .i_sdma_0_init_ht_0_axi_s_arcache       (sdma_0_to_center_init_ht_0_axi_arcache),
        .i_sdma_0_init_ht_0_axi_s_arid          (sdma_0_to_center_init_ht_0_axi_arid),
        .i_sdma_0_init_ht_0_axi_s_arlen         (sdma_0_to_center_init_ht_0_axi_arlen),
        .i_sdma_0_init_ht_0_axi_s_arlock        (sdma_0_to_center_init_ht_0_axi_arlock),
        .i_sdma_0_init_ht_0_axi_s_arprot        (sdma_0_to_center_init_ht_0_axi_arprot),
        .o_sdma_0_init_ht_0_axi_s_arready       (sdma_0_to_center_init_ht_0_axi_arready),
        .i_sdma_0_init_ht_0_axi_s_arsize        (sdma_0_to_center_init_ht_0_axi_arsize),
        .i_sdma_0_init_ht_0_axi_s_arvalid       (sdma_0_to_center_init_ht_0_axi_arvalid),
        .o_sdma_0_init_ht_0_axi_s_rdata         (sdma_0_to_center_init_ht_0_axi_rdata),
        .o_sdma_0_init_ht_0_axi_s_rid           (sdma_0_to_center_init_ht_0_axi_rid),
        .o_sdma_0_init_ht_0_axi_s_rlast         (sdma_0_to_center_init_ht_0_axi_rlast),
        .i_sdma_0_init_ht_0_axi_s_rready        (sdma_0_to_center_init_ht_0_axi_rready),
        .o_sdma_0_init_ht_0_axi_s_rresp         (sdma_0_to_center_init_ht_0_axi_rresp),
        .o_sdma_0_init_ht_0_axi_s_rvalid        (sdma_0_to_center_init_ht_0_axi_rvalid),
        .i_sdma_0_init_ht_0_axi_s_awaddr        (sdma_0_to_center_init_ht_0_axi_awaddr),
        .i_sdma_0_init_ht_0_axi_s_awburst       (sdma_0_to_center_init_ht_0_axi_awburst),
        .i_sdma_0_init_ht_0_axi_s_awcache       (sdma_0_to_center_init_ht_0_axi_awcache),
        .i_sdma_0_init_ht_0_axi_s_awid          (sdma_0_to_center_init_ht_0_axi_awid),
        .i_sdma_0_init_ht_0_axi_s_awlen         (sdma_0_to_center_init_ht_0_axi_awlen),
        .i_sdma_0_init_ht_0_axi_s_awlock        (sdma_0_to_center_init_ht_0_axi_awlock),
        .i_sdma_0_init_ht_0_axi_s_awprot        (sdma_0_to_center_init_ht_0_axi_awprot),
        .o_sdma_0_init_ht_0_axi_s_awready       (sdma_0_to_center_init_ht_0_axi_awready),
        .i_sdma_0_init_ht_0_axi_s_awsize        (sdma_0_to_center_init_ht_0_axi_awsize),
        .i_sdma_0_init_ht_0_axi_s_awvalid       (sdma_0_to_center_init_ht_0_axi_awvalid),
        .o_sdma_0_init_ht_0_axi_s_bid           (sdma_0_to_center_init_ht_0_axi_bid),
        .i_sdma_0_init_ht_0_axi_s_bready        (sdma_0_to_center_init_ht_0_axi_bready),
        .o_sdma_0_init_ht_0_axi_s_bresp         (sdma_0_to_center_init_ht_0_axi_bresp),
        .o_sdma_0_init_ht_0_axi_s_bvalid        (sdma_0_to_center_init_ht_0_axi_bvalid),
        .i_sdma_0_init_ht_0_axi_s_wdata         (sdma_0_to_center_init_ht_0_axi_wdata),
        .i_sdma_0_init_ht_0_axi_s_wlast         (sdma_0_to_center_init_ht_0_axi_wlast),
        .o_sdma_0_init_ht_0_axi_s_wready        (sdma_0_to_center_init_ht_0_axi_wready),
        .i_sdma_0_init_ht_0_axi_s_wstrb         (sdma_0_to_center_init_ht_0_axi_wstrb),
        .i_sdma_0_init_ht_0_axi_s_wvalid        (sdma_0_to_center_init_ht_0_axi_wvalid),
        .i_sdma_0_init_ht_1_axi_s_araddr        (sdma_0_to_center_init_ht_1_axi_araddr),
        .i_sdma_0_init_ht_1_axi_s_arburst       (sdma_0_to_center_init_ht_1_axi_arburst),
        .i_sdma_0_init_ht_1_axi_s_arcache       (sdma_0_to_center_init_ht_1_axi_arcache),
        .i_sdma_0_init_ht_1_axi_s_arid          (sdma_0_to_center_init_ht_1_axi_arid),
        .i_sdma_0_init_ht_1_axi_s_arlen         (sdma_0_to_center_init_ht_1_axi_arlen),
        .i_sdma_0_init_ht_1_axi_s_arlock        (sdma_0_to_center_init_ht_1_axi_arlock),
        .i_sdma_0_init_ht_1_axi_s_arprot        (sdma_0_to_center_init_ht_1_axi_arprot),
        .o_sdma_0_init_ht_1_axi_s_arready       (sdma_0_to_center_init_ht_1_axi_arready),
        .i_sdma_0_init_ht_1_axi_s_arsize        (sdma_0_to_center_init_ht_1_axi_arsize),
        .i_sdma_0_init_ht_1_axi_s_arvalid       (sdma_0_to_center_init_ht_1_axi_arvalid),
        .o_sdma_0_init_ht_1_axi_s_rdata         (sdma_0_to_center_init_ht_1_axi_rdata),
        .o_sdma_0_init_ht_1_axi_s_rid           (sdma_0_to_center_init_ht_1_axi_rid),
        .o_sdma_0_init_ht_1_axi_s_rlast         (sdma_0_to_center_init_ht_1_axi_rlast),
        .i_sdma_0_init_ht_1_axi_s_rready        (sdma_0_to_center_init_ht_1_axi_rready),
        .o_sdma_0_init_ht_1_axi_s_rresp         (sdma_0_to_center_init_ht_1_axi_rresp),
        .o_sdma_0_init_ht_1_axi_s_rvalid        (sdma_0_to_center_init_ht_1_axi_rvalid),
        .i_sdma_0_init_ht_1_axi_s_awaddr        (sdma_0_to_center_init_ht_1_axi_awaddr),
        .i_sdma_0_init_ht_1_axi_s_awburst       (sdma_0_to_center_init_ht_1_axi_awburst),
        .i_sdma_0_init_ht_1_axi_s_awcache       (sdma_0_to_center_init_ht_1_axi_awcache),
        .i_sdma_0_init_ht_1_axi_s_awid          (sdma_0_to_center_init_ht_1_axi_awid),
        .i_sdma_0_init_ht_1_axi_s_awlen         (sdma_0_to_center_init_ht_1_axi_awlen),
        .i_sdma_0_init_ht_1_axi_s_awlock        (sdma_0_to_center_init_ht_1_axi_awlock),
        .i_sdma_0_init_ht_1_axi_s_awprot        (sdma_0_to_center_init_ht_1_axi_awprot),
        .o_sdma_0_init_ht_1_axi_s_awready       (sdma_0_to_center_init_ht_1_axi_awready),
        .i_sdma_0_init_ht_1_axi_s_awsize        (sdma_0_to_center_init_ht_1_axi_awsize),
        .i_sdma_0_init_ht_1_axi_s_awvalid       (sdma_0_to_center_init_ht_1_axi_awvalid),
        .o_sdma_0_init_ht_1_axi_s_bid           (sdma_0_to_center_init_ht_1_axi_bid),
        .i_sdma_0_init_ht_1_axi_s_bready        (sdma_0_to_center_init_ht_1_axi_bready),
        .o_sdma_0_init_ht_1_axi_s_bresp         (sdma_0_to_center_init_ht_1_axi_bresp),
        .o_sdma_0_init_ht_1_axi_s_bvalid        (sdma_0_to_center_init_ht_1_axi_bvalid),
        .i_sdma_0_init_ht_1_axi_s_wdata         (sdma_0_to_center_init_ht_1_axi_wdata),
        .i_sdma_0_init_ht_1_axi_s_wlast         (sdma_0_to_center_init_ht_1_axi_wlast),
        .o_sdma_0_init_ht_1_axi_s_wready        (sdma_0_to_center_init_ht_1_axi_wready),
        .i_sdma_0_init_ht_1_axi_s_wstrb         (sdma_0_to_center_init_ht_1_axi_wstrb),
        .i_sdma_0_init_ht_1_axi_s_wvalid        (sdma_0_to_center_init_ht_1_axi_wvalid),
        .i_sdma_0_init_lt_axi_s_araddr          (sdma_0_to_center_init_lt_araddr),
        .i_sdma_0_init_lt_axi_s_arburst         (sdma_0_to_center_init_lt_arburst),
        .i_sdma_0_init_lt_axi_s_arcache         (sdma_0_to_center_init_lt_arcache),
        .i_sdma_0_init_lt_axi_s_arid            (sdma_0_to_center_init_lt_arid),
        .i_sdma_0_init_lt_axi_s_arlen           (sdma_0_to_center_init_lt_arlen),
        .i_sdma_0_init_lt_axi_s_arlock          (sdma_0_to_center_init_lt_arlock),
        .i_sdma_0_init_lt_axi_s_arprot          (sdma_0_to_center_init_lt_arprot),
        .i_sdma_0_init_lt_axi_s_arqos           (sdma_0_to_center_init_lt_arqos),
        .o_sdma_0_init_lt_axi_s_arready         (sdma_0_to_center_init_lt_arready),
        .i_sdma_0_init_lt_axi_s_arsize          (sdma_0_to_center_init_lt_arsize),
        .i_sdma_0_init_lt_axi_s_arvalid         (sdma_0_to_center_init_lt_arvalid),
        .i_sdma_0_init_lt_axi_s_awaddr          (sdma_0_to_center_init_lt_awaddr),
        .i_sdma_0_init_lt_axi_s_awburst         (sdma_0_to_center_init_lt_awburst),
        .i_sdma_0_init_lt_axi_s_awcache         (sdma_0_to_center_init_lt_awcache),
        .i_sdma_0_init_lt_axi_s_awid            (sdma_0_to_center_init_lt_awid),
        .i_sdma_0_init_lt_axi_s_awlen           (sdma_0_to_center_init_lt_awlen),
        .i_sdma_0_init_lt_axi_s_awlock          (sdma_0_to_center_init_lt_awlock),
        .i_sdma_0_init_lt_axi_s_awprot          (sdma_0_to_center_init_lt_awprot),
        .i_sdma_0_init_lt_axi_s_awqos           (sdma_0_to_center_init_lt_awqos),
        .o_sdma_0_init_lt_axi_s_awready         (sdma_0_to_center_init_lt_awready),
        .i_sdma_0_init_lt_axi_s_awsize          (sdma_0_to_center_init_lt_awsize),
        .i_sdma_0_init_lt_axi_s_awvalid         (sdma_0_to_center_init_lt_awvalid),
        .o_sdma_0_init_lt_axi_s_bid             (sdma_0_to_center_init_lt_bid),
        .i_sdma_0_init_lt_axi_s_bready          (sdma_0_to_center_init_lt_bready),
        .o_sdma_0_init_lt_axi_s_bresp           (sdma_0_to_center_init_lt_bresp),
        .o_sdma_0_init_lt_axi_s_bvalid          (sdma_0_to_center_init_lt_bvalid),
        .o_sdma_0_init_lt_axi_s_rdata           (sdma_0_to_center_init_lt_rdata),
        .o_sdma_0_init_lt_axi_s_rid             (sdma_0_to_center_init_lt_rid),
        .o_sdma_0_init_lt_axi_s_rlast           (sdma_0_to_center_init_lt_rlast),
        .i_sdma_0_init_lt_axi_s_rready          (sdma_0_to_center_init_lt_rready),
        .o_sdma_0_init_lt_axi_s_rresp           (sdma_0_to_center_init_lt_rresp),
        .o_sdma_0_init_lt_axi_s_rvalid          (sdma_0_to_center_init_lt_rvalid),
        .i_sdma_0_init_lt_axi_s_wdata           (sdma_0_to_center_init_lt_wdata),
        .i_sdma_0_init_lt_axi_s_wlast           (sdma_0_to_center_init_lt_wlast),
        .o_sdma_0_init_lt_axi_s_wready          (sdma_0_to_center_init_lt_wready),
        .i_sdma_0_init_lt_axi_s_wstrb           (sdma_0_to_center_init_lt_wstrb),
        .i_sdma_0_init_lt_axi_s_wvalid          (sdma_0_to_center_init_lt_wvalid),
        .o_sdma_0_pwr_idle_val                  (center_to_sdma_0_noc_async_idle_val),
        .o_sdma_0_pwr_idle_ack                  (center_to_sdma_0_noc_async_idle_ack),
        .i_sdma_0_pwr_idle_req                  (center_to_sdma_0_noc_async_idle_req),
        .i_sdma_0_rst_n                         (center_to_sdma_0_noc_rst_n),
        .o_sdma_0_targ_lt_axi_m_araddr          (center_to_sdma_0_targ_lt_axi_araddr),
        .o_sdma_0_targ_lt_axi_m_arburst         (center_to_sdma_0_targ_lt_axi_arburst),
        .o_sdma_0_targ_lt_axi_m_arcache         (center_to_sdma_0_targ_lt_axi_arcache),
        .o_sdma_0_targ_lt_axi_m_arid            (center_to_sdma_0_targ_lt_axi_arid),
        .o_sdma_0_targ_lt_axi_m_arlen           (center_to_sdma_0_targ_lt_axi_arlen),
        .o_sdma_0_targ_lt_axi_m_arlock          (center_to_sdma_0_targ_lt_axi_arlock),
        .o_sdma_0_targ_lt_axi_m_arprot          (center_to_sdma_0_targ_lt_axi_arprot),
        .o_sdma_0_targ_lt_axi_m_arqos           ( ),  // TODO(psarras; bronze; confirm this is unused)
        .i_sdma_0_targ_lt_axi_m_arready         (center_to_sdma_0_targ_lt_axi_arready),
        .o_sdma_0_targ_lt_axi_m_arsize          (center_to_sdma_0_targ_lt_axi_arsize),
        .o_sdma_0_targ_lt_axi_m_arvalid         (center_to_sdma_0_targ_lt_axi_arvalid),
        .o_sdma_0_targ_lt_axi_m_awaddr          (center_to_sdma_0_targ_lt_axi_awaddr),
        .o_sdma_0_targ_lt_axi_m_awburst         (center_to_sdma_0_targ_lt_axi_awburst),
        .o_sdma_0_targ_lt_axi_m_awcache         (center_to_sdma_0_targ_lt_axi_awcache),
        .o_sdma_0_targ_lt_axi_m_awid            (center_to_sdma_0_targ_lt_axi_awid),
        .o_sdma_0_targ_lt_axi_m_awlen           (center_to_sdma_0_targ_lt_axi_awlen),
        .o_sdma_0_targ_lt_axi_m_awlock          (center_to_sdma_0_targ_lt_axi_awlock),
        .o_sdma_0_targ_lt_axi_m_awprot          (center_to_sdma_0_targ_lt_axi_awprot),
        .o_sdma_0_targ_lt_axi_m_awqos           ( ), // TODO(psarras; bronze; confirm this is unused)
        .i_sdma_0_targ_lt_axi_m_awready         (center_to_sdma_0_targ_lt_axi_awready),
        .o_sdma_0_targ_lt_axi_m_awsize          (center_to_sdma_0_targ_lt_axi_awsize),
        .o_sdma_0_targ_lt_axi_m_awvalid         (center_to_sdma_0_targ_lt_axi_awvalid),
        .i_sdma_0_targ_lt_axi_m_bid             (center_to_sdma_0_targ_lt_axi_bid),
        .o_sdma_0_targ_lt_axi_m_bready          (center_to_sdma_0_targ_lt_axi_bready),
        .i_sdma_0_targ_lt_axi_m_bresp           (center_to_sdma_0_targ_lt_axi_bresp),
        .i_sdma_0_targ_lt_axi_m_bvalid          (center_to_sdma_0_targ_lt_axi_bvalid),
        .i_sdma_0_targ_lt_axi_m_rdata           (center_to_sdma_0_targ_lt_axi_rdata),
        .i_sdma_0_targ_lt_axi_m_rid             (center_to_sdma_0_targ_lt_axi_rid),
        .i_sdma_0_targ_lt_axi_m_rlast           (center_to_sdma_0_targ_lt_axi_rlast),
        .o_sdma_0_targ_lt_axi_m_rready          (center_to_sdma_0_targ_lt_axi_rready),
        .i_sdma_0_targ_lt_axi_m_rresp           (center_to_sdma_0_targ_lt_axi_rresp),
        .i_sdma_0_targ_lt_axi_m_rvalid          (center_to_sdma_0_targ_lt_axi_rvalid),
        .o_sdma_0_targ_lt_axi_m_wdata           (center_to_sdma_0_targ_lt_axi_wdata),
        .o_sdma_0_targ_lt_axi_m_wlast           (center_to_sdma_0_targ_lt_axi_wlast),
        .i_sdma_0_targ_lt_axi_m_wready          (center_to_sdma_0_targ_lt_axi_wready),
        .o_sdma_0_targ_lt_axi_m_wstrb           (center_to_sdma_0_targ_lt_axi_wstrb),
        .o_sdma_0_targ_lt_axi_m_wvalid          (center_to_sdma_0_targ_lt_axi_wvalid),
        .o_sdma_0_targ_syscfg_apb_m_paddr       (center_to_sdma_0_cfg_apb4_paddr),
        .o_sdma_0_targ_syscfg_apb_m_penable     (center_to_sdma_0_cfg_apb4_penable),
        .o_sdma_0_targ_syscfg_apb_m_pprot       (center_to_sdma_0_cfg_apb4_pprot),
        .i_sdma_0_targ_syscfg_apb_m_prdata      (center_to_sdma_0_cfg_apb4_prdata),
        .i_sdma_0_targ_syscfg_apb_m_pready      (center_to_sdma_0_cfg_apb4_pready),
        .o_sdma_0_targ_syscfg_apb_m_psel        (center_to_sdma_0_cfg_apb4_psel),
        .i_sdma_0_targ_syscfg_apb_m_pslverr     (center_to_sdma_0_cfg_apb4_pslverr),
        .o_sdma_0_targ_syscfg_apb_m_pstrb       (center_to_sdma_0_cfg_apb4_pstrb),
        .o_sdma_0_targ_syscfg_apb_m_pwdata      (center_to_sdma_0_cfg_apb4_pwdata),
        .o_sdma_0_targ_syscfg_apb_m_pwrite      (center_to_sdma_0_cfg_apb4_pwrite),

        .i_sdma_1_aon_clk                       (i_ref_clk),
        .i_sdma_1_aon_rst_n                     (i_sdma_1_ao_rst_n),
        .i_sdma_1_clk                           (i_sdma_1_clk),
        .i_sdma_1_clken                         (center_to_sdma_1_noc_clken),
        .i_sdma_1_init_ht_0_axi_s_araddr        (sdma_1_to_center_init_ht_0_axi_araddr),
        .i_sdma_1_init_ht_0_axi_s_arburst       (sdma_1_to_center_init_ht_0_axi_arburst),
        .i_sdma_1_init_ht_0_axi_s_arcache       (sdma_1_to_center_init_ht_0_axi_arcache),
        .i_sdma_1_init_ht_0_axi_s_arid          (sdma_1_to_center_init_ht_0_axi_arid),
        .i_sdma_1_init_ht_0_axi_s_arlen         (sdma_1_to_center_init_ht_0_axi_arlen),
        .i_sdma_1_init_ht_0_axi_s_arlock        (sdma_1_to_center_init_ht_0_axi_arlock),
        .i_sdma_1_init_ht_0_axi_s_arprot        (sdma_1_to_center_init_ht_0_axi_arprot),
        .o_sdma_1_init_ht_0_axi_s_arready       (sdma_1_to_center_init_ht_0_axi_arready),
        .i_sdma_1_init_ht_0_axi_s_arsize        (sdma_1_to_center_init_ht_0_axi_arsize),
        .i_sdma_1_init_ht_0_axi_s_arvalid       (sdma_1_to_center_init_ht_0_axi_arvalid),
        .o_sdma_1_init_ht_0_axi_s_rdata         (sdma_1_to_center_init_ht_0_axi_rdata),
        .o_sdma_1_init_ht_0_axi_s_rid           (sdma_1_to_center_init_ht_0_axi_rid),
        .o_sdma_1_init_ht_0_axi_s_rlast         (sdma_1_to_center_init_ht_0_axi_rlast),
        .i_sdma_1_init_ht_0_axi_s_rready        (sdma_1_to_center_init_ht_0_axi_rready),
        .o_sdma_1_init_ht_0_axi_s_rresp         (sdma_1_to_center_init_ht_0_axi_rresp),
        .o_sdma_1_init_ht_0_axi_s_rvalid        (sdma_1_to_center_init_ht_0_axi_rvalid),
        .i_sdma_1_init_ht_0_axi_s_awaddr        (sdma_1_to_center_init_ht_0_axi_awaddr),
        .i_sdma_1_init_ht_0_axi_s_awburst       (sdma_1_to_center_init_ht_0_axi_awburst),
        .i_sdma_1_init_ht_0_axi_s_awcache       (sdma_1_to_center_init_ht_0_axi_awcache),
        .i_sdma_1_init_ht_0_axi_s_awid          (sdma_1_to_center_init_ht_0_axi_awid),
        .i_sdma_1_init_ht_0_axi_s_awlen         (sdma_1_to_center_init_ht_0_axi_awlen),
        .i_sdma_1_init_ht_0_axi_s_awlock        (sdma_1_to_center_init_ht_0_axi_awlock),
        .i_sdma_1_init_ht_0_axi_s_awprot        (sdma_1_to_center_init_ht_0_axi_awprot),
        .o_sdma_1_init_ht_0_axi_s_awready       (sdma_1_to_center_init_ht_0_axi_awready),
        .i_sdma_1_init_ht_0_axi_s_awsize        (sdma_1_to_center_init_ht_0_axi_awsize),
        .i_sdma_1_init_ht_0_axi_s_awvalid       (sdma_1_to_center_init_ht_0_axi_awvalid),
        .o_sdma_1_init_ht_0_axi_s_bid           (sdma_1_to_center_init_ht_0_axi_bid),
        .i_sdma_1_init_ht_0_axi_s_bready        (sdma_1_to_center_init_ht_0_axi_bready),
        .o_sdma_1_init_ht_0_axi_s_bresp         (sdma_1_to_center_init_ht_0_axi_bresp),
        .o_sdma_1_init_ht_0_axi_s_bvalid        (sdma_1_to_center_init_ht_0_axi_bvalid),
        .i_sdma_1_init_ht_0_axi_s_wdata         (sdma_1_to_center_init_ht_0_axi_wdata),
        .i_sdma_1_init_ht_0_axi_s_wlast         (sdma_1_to_center_init_ht_0_axi_wlast),
        .o_sdma_1_init_ht_0_axi_s_wready        (sdma_1_to_center_init_ht_0_axi_wready),
        .i_sdma_1_init_ht_0_axi_s_wstrb         (sdma_1_to_center_init_ht_0_axi_wstrb),
        .i_sdma_1_init_ht_0_axi_s_wvalid        (sdma_1_to_center_init_ht_0_axi_wvalid),
        .i_sdma_1_init_ht_1_axi_s_araddr        (sdma_1_to_center_init_ht_1_axi_araddr),
        .i_sdma_1_init_ht_1_axi_s_arburst       (sdma_1_to_center_init_ht_1_axi_arburst),
        .i_sdma_1_init_ht_1_axi_s_arcache       (sdma_1_to_center_init_ht_1_axi_arcache),
        .i_sdma_1_init_ht_1_axi_s_arid          (sdma_1_to_center_init_ht_1_axi_arid),
        .i_sdma_1_init_ht_1_axi_s_arlen         (sdma_1_to_center_init_ht_1_axi_arlen),
        .i_sdma_1_init_ht_1_axi_s_arlock        (sdma_1_to_center_init_ht_1_axi_arlock),
        .i_sdma_1_init_ht_1_axi_s_arprot        (sdma_1_to_center_init_ht_1_axi_arprot),
        .o_sdma_1_init_ht_1_axi_s_arready       (sdma_1_to_center_init_ht_1_axi_arready),
        .i_sdma_1_init_ht_1_axi_s_arsize        (sdma_1_to_center_init_ht_1_axi_arsize),
        .i_sdma_1_init_ht_1_axi_s_arvalid       (sdma_1_to_center_init_ht_1_axi_arvalid),
        .o_sdma_1_init_ht_1_axi_s_rdata         (sdma_1_to_center_init_ht_1_axi_rdata),
        .o_sdma_1_init_ht_1_axi_s_rid           (sdma_1_to_center_init_ht_1_axi_rid),
        .o_sdma_1_init_ht_1_axi_s_rlast         (sdma_1_to_center_init_ht_1_axi_rlast),
        .i_sdma_1_init_ht_1_axi_s_rready        (sdma_1_to_center_init_ht_1_axi_rready),
        .o_sdma_1_init_ht_1_axi_s_rresp         (sdma_1_to_center_init_ht_1_axi_rresp),
        .o_sdma_1_init_ht_1_axi_s_rvalid        (sdma_1_to_center_init_ht_1_axi_rvalid),
        .i_sdma_1_init_ht_1_axi_s_awaddr        (sdma_1_to_center_init_ht_1_axi_awaddr),
        .i_sdma_1_init_ht_1_axi_s_awburst       (sdma_1_to_center_init_ht_1_axi_awburst),
        .i_sdma_1_init_ht_1_axi_s_awcache       (sdma_1_to_center_init_ht_1_axi_awcache),
        .i_sdma_1_init_ht_1_axi_s_awid          (sdma_1_to_center_init_ht_1_axi_awid),
        .i_sdma_1_init_ht_1_axi_s_awlen         (sdma_1_to_center_init_ht_1_axi_awlen),
        .i_sdma_1_init_ht_1_axi_s_awlock        (sdma_1_to_center_init_ht_1_axi_awlock),
        .i_sdma_1_init_ht_1_axi_s_awprot        (sdma_1_to_center_init_ht_1_axi_awprot),
        .o_sdma_1_init_ht_1_axi_s_awready       (sdma_1_to_center_init_ht_1_axi_awready),
        .i_sdma_1_init_ht_1_axi_s_awsize        (sdma_1_to_center_init_ht_1_axi_awsize),
        .i_sdma_1_init_ht_1_axi_s_awvalid       (sdma_1_to_center_init_ht_1_axi_awvalid),
        .o_sdma_1_init_ht_1_axi_s_bid           (sdma_1_to_center_init_ht_1_axi_bid),
        .i_sdma_1_init_ht_1_axi_s_bready        (sdma_1_to_center_init_ht_1_axi_bready),
        .o_sdma_1_init_ht_1_axi_s_bresp         (sdma_1_to_center_init_ht_1_axi_bresp),
        .o_sdma_1_init_ht_1_axi_s_bvalid        (sdma_1_to_center_init_ht_1_axi_bvalid),
        .i_sdma_1_init_ht_1_axi_s_wdata         (sdma_1_to_center_init_ht_1_axi_wdata),
        .i_sdma_1_init_ht_1_axi_s_wlast         (sdma_1_to_center_init_ht_1_axi_wlast),
        .o_sdma_1_init_ht_1_axi_s_wready        (sdma_1_to_center_init_ht_1_axi_wready),
        .i_sdma_1_init_ht_1_axi_s_wstrb         (sdma_1_to_center_init_ht_1_axi_wstrb),
        .i_sdma_1_init_ht_1_axi_s_wvalid        (sdma_1_to_center_init_ht_1_axi_wvalid),
        .i_sdma_1_init_lt_axi_s_araddr          (sdma_1_to_center_init_lt_araddr),
        .i_sdma_1_init_lt_axi_s_arburst         (sdma_1_to_center_init_lt_arburst),
        .i_sdma_1_init_lt_axi_s_arcache         (sdma_1_to_center_init_lt_arcache),
        .i_sdma_1_init_lt_axi_s_arid            (sdma_1_to_center_init_lt_arid),
        .i_sdma_1_init_lt_axi_s_arlen           (sdma_1_to_center_init_lt_arlen),
        .i_sdma_1_init_lt_axi_s_arlock          (sdma_1_to_center_init_lt_arlock),
        .i_sdma_1_init_lt_axi_s_arprot          (sdma_1_to_center_init_lt_arprot),
        .i_sdma_1_init_lt_axi_s_arqos           (sdma_1_to_center_init_lt_arqos),
        .o_sdma_1_init_lt_axi_s_arready         (sdma_1_to_center_init_lt_arready),
        .i_sdma_1_init_lt_axi_s_arsize          (sdma_1_to_center_init_lt_arsize),
        .i_sdma_1_init_lt_axi_s_arvalid         (sdma_1_to_center_init_lt_arvalid),
        .i_sdma_1_init_lt_axi_s_awaddr          (sdma_1_to_center_init_lt_awaddr),
        .i_sdma_1_init_lt_axi_s_awburst         (sdma_1_to_center_init_lt_awburst),
        .i_sdma_1_init_lt_axi_s_awcache         (sdma_1_to_center_init_lt_awcache),
        .i_sdma_1_init_lt_axi_s_awid            (sdma_1_to_center_init_lt_awid),
        .i_sdma_1_init_lt_axi_s_awlen           (sdma_1_to_center_init_lt_awlen),
        .i_sdma_1_init_lt_axi_s_awlock          (sdma_1_to_center_init_lt_awlock),
        .i_sdma_1_init_lt_axi_s_awprot          (sdma_1_to_center_init_lt_awprot),
        .i_sdma_1_init_lt_axi_s_awqos           (sdma_1_to_center_init_lt_awqos),
        .o_sdma_1_init_lt_axi_s_awready         (sdma_1_to_center_init_lt_awready),
        .i_sdma_1_init_lt_axi_s_awsize          (sdma_1_to_center_init_lt_awsize),
        .i_sdma_1_init_lt_axi_s_awvalid         (sdma_1_to_center_init_lt_awvalid),
        .o_sdma_1_init_lt_axi_s_bid             (sdma_1_to_center_init_lt_bid),
        .i_sdma_1_init_lt_axi_s_bready          (sdma_1_to_center_init_lt_bready),
        .o_sdma_1_init_lt_axi_s_bresp           (sdma_1_to_center_init_lt_bresp),
        .o_sdma_1_init_lt_axi_s_bvalid          (sdma_1_to_center_init_lt_bvalid),
        .o_sdma_1_init_lt_axi_s_rdata           (sdma_1_to_center_init_lt_rdata),
        .o_sdma_1_init_lt_axi_s_rid             (sdma_1_to_center_init_lt_rid),
        .o_sdma_1_init_lt_axi_s_rlast           (sdma_1_to_center_init_lt_rlast),
        .i_sdma_1_init_lt_axi_s_rready          (sdma_1_to_center_init_lt_rready),
        .o_sdma_1_init_lt_axi_s_rresp           (sdma_1_to_center_init_lt_rresp),
        .o_sdma_1_init_lt_axi_s_rvalid          (sdma_1_to_center_init_lt_rvalid),
        .i_sdma_1_init_lt_axi_s_wdata           (sdma_1_to_center_init_lt_wdata),
        .i_sdma_1_init_lt_axi_s_wlast           (sdma_1_to_center_init_lt_wlast),
        .o_sdma_1_init_lt_axi_s_wready          (sdma_1_to_center_init_lt_wready),
        .i_sdma_1_init_lt_axi_s_wstrb           (sdma_1_to_center_init_lt_wstrb),
        .i_sdma_1_init_lt_axi_s_wvalid          (sdma_1_to_center_init_lt_wvalid),
        .o_sdma_1_pwr_idle_val                  (center_to_sdma_1_noc_async_idle_val),
        .o_sdma_1_pwr_idle_ack                  (center_to_sdma_1_noc_async_idle_ack),
        .i_sdma_1_pwr_idle_req                  (center_to_sdma_1_noc_async_idle_req),
        .i_sdma_1_rst_n                         (center_to_sdma_1_noc_rst_n),
        .o_sdma_1_targ_lt_axi_m_araddr          (center_to_sdma_1_targ_lt_axi_araddr),
        .o_sdma_1_targ_lt_axi_m_arburst         (center_to_sdma_1_targ_lt_axi_arburst),
        .o_sdma_1_targ_lt_axi_m_arcache         (center_to_sdma_1_targ_lt_axi_arcache),
        .o_sdma_1_targ_lt_axi_m_arid            (center_to_sdma_1_targ_lt_axi_arid),
        .o_sdma_1_targ_lt_axi_m_arlen           (center_to_sdma_1_targ_lt_axi_arlen),
        .o_sdma_1_targ_lt_axi_m_arlock          (center_to_sdma_1_targ_lt_axi_arlock),
        .o_sdma_1_targ_lt_axi_m_arprot          (center_to_sdma_1_targ_lt_axi_arprot),
        .o_sdma_1_targ_lt_axi_m_arqos           ( ), // TODO(psarras; bronze; confirm this is unused)
        .i_sdma_1_targ_lt_axi_m_arready         (center_to_sdma_1_targ_lt_axi_arready),
        .o_sdma_1_targ_lt_axi_m_arsize          (center_to_sdma_1_targ_lt_axi_arsize),
        .o_sdma_1_targ_lt_axi_m_arvalid         (center_to_sdma_1_targ_lt_axi_arvalid),
        .o_sdma_1_targ_lt_axi_m_awaddr          (center_to_sdma_1_targ_lt_axi_awaddr),
        .o_sdma_1_targ_lt_axi_m_awburst         (center_to_sdma_1_targ_lt_axi_awburst),
        .o_sdma_1_targ_lt_axi_m_awcache         (center_to_sdma_1_targ_lt_axi_awcache),
        .o_sdma_1_targ_lt_axi_m_awid            (center_to_sdma_1_targ_lt_axi_awid),
        .o_sdma_1_targ_lt_axi_m_awlen           (center_to_sdma_1_targ_lt_axi_awlen),
        .o_sdma_1_targ_lt_axi_m_awlock          (center_to_sdma_1_targ_lt_axi_awlock),
        .o_sdma_1_targ_lt_axi_m_awprot          (center_to_sdma_1_targ_lt_axi_awprot),
        .o_sdma_1_targ_lt_axi_m_awqos           ( ),  // TODO(psarras; bronze; confirm this is unused)
        .i_sdma_1_targ_lt_axi_m_awready         (center_to_sdma_1_targ_lt_axi_awready),
        .o_sdma_1_targ_lt_axi_m_awsize          (center_to_sdma_1_targ_lt_axi_awsize),
        .o_sdma_1_targ_lt_axi_m_awvalid         (center_to_sdma_1_targ_lt_axi_awvalid),
        .i_sdma_1_targ_lt_axi_m_bid             (center_to_sdma_1_targ_lt_axi_bid),
        .o_sdma_1_targ_lt_axi_m_bready          (center_to_sdma_1_targ_lt_axi_bready),
        .i_sdma_1_targ_lt_axi_m_bresp           (center_to_sdma_1_targ_lt_axi_bresp),
        .i_sdma_1_targ_lt_axi_m_bvalid          (center_to_sdma_1_targ_lt_axi_bvalid),
        .i_sdma_1_targ_lt_axi_m_rdata           (center_to_sdma_1_targ_lt_axi_rdata),
        .i_sdma_1_targ_lt_axi_m_rid             (center_to_sdma_1_targ_lt_axi_rid),
        .i_sdma_1_targ_lt_axi_m_rlast           (center_to_sdma_1_targ_lt_axi_rlast),
        .o_sdma_1_targ_lt_axi_m_rready          (center_to_sdma_1_targ_lt_axi_rready),
        .i_sdma_1_targ_lt_axi_m_rresp           (center_to_sdma_1_targ_lt_axi_rresp),
        .i_sdma_1_targ_lt_axi_m_rvalid          (center_to_sdma_1_targ_lt_axi_rvalid),
        .o_sdma_1_targ_lt_axi_m_wdata           (center_to_sdma_1_targ_lt_axi_wdata),
        .o_sdma_1_targ_lt_axi_m_wlast           (center_to_sdma_1_targ_lt_axi_wlast),
        .i_sdma_1_targ_lt_axi_m_wready          (center_to_sdma_1_targ_lt_axi_wready),
        .o_sdma_1_targ_lt_axi_m_wstrb           (center_to_sdma_1_targ_lt_axi_wstrb),
        .o_sdma_1_targ_lt_axi_m_wvalid          (center_to_sdma_1_targ_lt_axi_wvalid),
        .o_sdma_1_targ_syscfg_apb_m_paddr       (center_to_sdma_1_cfg_apb4_paddr),
        .o_sdma_1_targ_syscfg_apb_m_penable     (center_to_sdma_1_cfg_apb4_penable),
        .o_sdma_1_targ_syscfg_apb_m_pprot       (center_to_sdma_1_cfg_apb4_pprot),
        .i_sdma_1_targ_syscfg_apb_m_prdata      (center_to_sdma_1_cfg_apb4_prdata),
        .i_sdma_1_targ_syscfg_apb_m_pready      (center_to_sdma_1_cfg_apb4_pready),
        .o_sdma_1_targ_syscfg_apb_m_psel        (center_to_sdma_1_cfg_apb4_psel),
        .i_sdma_1_targ_syscfg_apb_m_pslverr     (center_to_sdma_1_cfg_apb4_pslverr),
        .o_sdma_1_targ_syscfg_apb_m_pstrb       (center_to_sdma_1_cfg_apb4_pstrb),
        .o_sdma_1_targ_syscfg_apb_m_pwdata      (center_to_sdma_1_cfg_apb4_pwdata),
        .o_sdma_1_targ_syscfg_apb_m_pwrite      (center_to_sdma_1_cfg_apb4_pwrite),

        .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld(dp_lnk_cross_center_to_east_512_0_egr_wr_req_to_lnk_cross_center_to_east_512_0_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld(dp_lnk_cross_center_to_east_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_0_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld(dp_lnk_cross_center_to_east_512_1_egr_wr_req_to_lnk_cross_center_to_east_512_1_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld(dp_lnk_cross_center_to_east_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_east_512_1_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld(dp_lnk_cross_center_to_east_512_2_egr_rd_req_to_lnk_cross_center_to_east_512_2_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld(dp_lnk_cross_center_to_east_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_2_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld(dp_lnk_cross_center_to_east_512_3_egr_rd_req_to_lnk_cross_center_to_east_512_3_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld(dp_lnk_cross_center_to_east_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_east_512_3_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_data),
        .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_head),
        .i_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_rdy),
        .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_tail),
        .o_dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld(dp_lnk_cross_center_to_east_64_egr_req_to_lnk_cross_center_to_east_64_ingr_req_vld),
        .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_data),
        .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_head),
        .o_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_tail),
        .i_dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld(dp_lnk_cross_center_to_east_64_ingr_req_resp_to_lnk_cross_center_to_east_64_egr_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_0_egr_wr_req_to_lnk_cross_center_to_north_512_0_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_0_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_1_egr_wr_req_to_lnk_cross_center_to_north_512_1_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_1_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_2_egr_rd_req_to_lnk_cross_center_to_north_512_2_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_2_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_3_egr_rd_req_to_lnk_cross_center_to_north_512_3_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_3_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_3_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_4_egr_rd_req_to_lnk_cross_center_to_north_512_4_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_4_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_5_egr_rd_req_to_lnk_cross_center_to_north_512_5_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_5_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_5_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_6_egr_wr_req_to_lnk_cross_center_to_north_512_6_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_6_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_6_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_7_egr_wr_req_to_lnk_cross_center_to_north_512_7_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_7_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_7_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_8_egr_wr_req_to_lnk_cross_center_to_north_512_8_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_8_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_9_egr_rd_req_to_lnk_cross_center_to_north_512_9_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_9_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld(dp_lnk_cross_center_to_north_512_a_egr_wr_req_to_lnk_cross_center_to_north_512_a_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld(dp_lnk_cross_center_to_north_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_north_512_a_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld(dp_lnk_cross_center_to_north_512_b_egr_rd_req_to_lnk_cross_center_to_north_512_b_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld(dp_lnk_cross_center_to_north_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_north_512_b_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_data),
        .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_head),
        .i_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_rdy),
        .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_tail),
        .o_dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld(dp_lnk_cross_center_to_north_64_egr_req_to_lnk_cross_center_to_north_64_ingr_req_vld),
        .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_data),
        .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_head),
        .o_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_tail),
        .i_dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld(dp_lnk_cross_center_to_north_64_ingr_req_resp_to_lnk_cross_center_to_north_64_egr_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_0_egr_wr_req_to_lnk_cross_center_to_south_512_0_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_0_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_0_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_1_egr_wr_req_to_lnk_cross_center_to_south_512_1_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_1_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_1_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_2_egr_rd_req_to_lnk_cross_center_to_south_512_2_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_2_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_2_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_3_egr_wr_req_to_lnk_cross_center_to_south_512_3_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_3_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_3_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_4_egr_rd_req_to_lnk_cross_center_to_south_512_4_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_4_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_4_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_5_egr_wr_req_to_lnk_cross_center_to_south_512_5_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_5_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_5_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_6_egr_rd_req_to_lnk_cross_center_to_south_512_6_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_6_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_6_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_7_egr_rd_req_to_lnk_cross_center_to_south_512_7_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_7_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_7_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_8_egr_wr_req_to_lnk_cross_center_to_south_512_8_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_8_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_8_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_9_egr_rd_req_to_lnk_cross_center_to_south_512_9_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_9_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_9_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_data),
        .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_head),
        .i_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_tail),
        .o_dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld(dp_lnk_cross_center_to_south_512_a_egr_wr_req_to_lnk_cross_center_to_south_512_a_ingr_wr_req_vld),
        .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld(dp_lnk_cross_center_to_south_512_a_ingr_wr_req_resp_to_lnk_cross_center_to_south_512_a_egr_wr_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_data),
        .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_head),
        .i_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_rdy),
        .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_tail),
        .o_dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld(dp_lnk_cross_center_to_south_512_b_egr_rd_req_to_lnk_cross_center_to_south_512_b_ingr_rd_req_vld),
        .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_data),
        .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_head),
        .o_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld(dp_lnk_cross_center_to_south_512_b_ingr_rd_req_resp_to_lnk_cross_center_to_south_512_b_egr_rd_req_resp_vld),
        .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_data),
        .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_head),
        .i_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_rdy),
        .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_tail),
        .o_dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld(dp_lnk_cross_center_to_south_64_egr_req_to_lnk_cross_center_to_south_64_ingr_req_vld),
        .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_data),
        .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_head),
        .o_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_rdy),
        .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_tail),
        .i_dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld(dp_lnk_cross_center_to_south_64_ingr_req_resp_to_lnk_cross_center_to_south_64_egr_req_resp_vld),
        .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_data),
        .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_head),
        .o_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_rdy),
        .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_tail),
        .i_dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld(dp_lnk_cross_center_to_west_32_ingr_resp_to_lnk_cross_center_to_west_64_egr_resp_vld),
        .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_data),
        .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_head),
        .i_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_rdy),
        .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_tail),
        .o_dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld(dp_lnk_cross_center_to_west_512_0_egr_to_lnk_cross_center_to_west_512_0_ingr_vld),
        .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_data),
        .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_head),
        .o_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_rdy),
        .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_tail),
        .i_dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld(dp_lnk_cross_center_to_west_512_0_ingr_resp_to_lnk_cross_center_to_west_512_0_egr_resp_vld),
        .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_data),
        .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_head),
        .i_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_rdy),
        .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_tail),
        .o_dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld(dp_lnk_cross_center_to_west_512_1_egr_to_lnk_cross_center_to_west_512_1_ingr_vld),
        .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_data),
        .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_head),
        .o_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_rdy),
        .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_tail),
        .i_dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld(dp_lnk_cross_center_to_west_512_1_ingr_resp_to_lnk_cross_center_to_west_512_1_egr_resp_vld),
        .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_data),
        .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_head),
        .i_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_rdy),
        .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_tail),
        .o_dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld(dp_lnk_cross_center_to_west_512_2_egr_to_lnk_cross_center_to_west_512_2_ingr_vld),
        .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_data),
        .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_head),
        .o_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_rdy),
        .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_tail),
        .i_dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld(dp_lnk_cross_center_to_west_512_2_ingr_resp_to_lnk_cross_center_to_west_512_2_egr_resp_vld),
        .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_data),
        .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_head),
        .i_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_rdy),
        .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_tail),
        .o_dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld(dp_lnk_cross_center_to_west_512_3_egr_to_lnk_cross_center_to_west_512_3_ingr_vld),
        .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_data),
        .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_head),
        .o_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_rdy),
        .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_tail),
        .i_dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld(dp_lnk_cross_center_to_west_512_3_ingr_resp_to_lnk_cross_center_to_west_512_3_egr_resp_vld),
        .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_data),
        .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_head),
        .i_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_rdy),
        .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_tail),
        .o_dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld(dp_lnk_cross_center_to_west_64_egr_to_lnk_cross_center_to_west_32_ingr_vld),
        .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_data),
        .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_head),
        .o_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_rdy),
        .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_tail),
        .i_dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld(dp_lnk_cross_east_to_center_512_0_egr_wr_req_to_lnk_cross_east_to_center_512_0_ingr_wr_req_vld),
        .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_data),
        .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_head),
        .i_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld(dp_lnk_cross_east_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_east_to_center_512_0_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_data),
        .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_head),
        .o_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_rdy),
        .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_tail),
        .i_dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld(dp_lnk_cross_east_to_center_512_1_egr_rd_req_to_lnk_cross_east_to_center_512_1_ingr_rd_req_vld),
        .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_data),
        .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_head),
        .i_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld(dp_lnk_cross_east_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_east_to_center_512_1_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_data),
        .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_head),
        .o_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_rdy),
        .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_tail),
        .i_dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld(dp_lnk_cross_east_to_center_64_egr_req_to_lnk_cross_east_to_center_64_ingr_req_vld),
        .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_data),
        .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_head),
        .i_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_tail),
        .o_dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld(dp_lnk_cross_east_to_center_64_ingr_req_resp_to_lnk_cross_east_to_center_64_egr_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_data),
        .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_head),
        .o_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_tail),
        .i_dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_0_egr_wr_req_to_lnk_cross_north_to_center_512_0_ingr_wr_req_vld),
        .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_0_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_0_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_data),
        .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_head),
        .o_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_tail),
        .i_dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_1_egr_rd_req_to_lnk_cross_north_to_center_512_1_ingr_rd_req_vld),
        .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_1_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_1_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_data),
        .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_head),
        .o_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_tail),
        .i_dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_2_egr_rd_req_to_lnk_cross_north_to_center_512_2_ingr_rd_req_vld),
        .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_2_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_2_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_data),
        .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_head),
        .o_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_tail),
        .i_dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_3_egr_rd_req_to_lnk_cross_north_to_center_512_3_ingr_rd_req_vld),
        .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_3_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_data),
        .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_head),
        .o_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_tail),
        .i_dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_4_egr_rd_req_to_lnk_cross_north_to_center_512_4_ingr_rd_req_vld),
        .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_4_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_data),
        .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_head),
        .o_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_tail),
        .i_dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_5_egr_rd_req_to_lnk_cross_north_to_center_512_5_ingr_rd_req_vld),
        .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_5_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_5_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_data),
        .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_head),
        .o_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_tail),
        .i_dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_6_egr_wr_req_to_lnk_cross_north_to_center_512_6_ingr_wr_req_vld),
        .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_6_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_data),
        .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_head),
        .o_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_tail),
        .i_dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_7_egr_wr_req_to_lnk_cross_north_to_center_512_7_ingr_wr_req_vld),
        .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_7_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_data),
        .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_head),
        .o_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_tail),
        .i_dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_8_egr_wr_req_to_lnk_cross_north_to_center_512_8_ingr_wr_req_vld),
        .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_8_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_8_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_data),
        .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_head),
        .o_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_tail),
        .i_dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_9_egr_wr_req_to_lnk_cross_north_to_center_512_9_ingr_wr_req_vld),
        .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_9_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_9_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_data),
        .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_head),
        .o_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_tail),
        .i_dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld(dp_lnk_cross_north_to_center_512_a_egr_wr_req_to_lnk_cross_north_to_center_512_a_ingr_wr_req_vld),
        .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld(dp_lnk_cross_north_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_north_to_center_512_a_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_data),
        .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_head),
        .o_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_rdy),
        .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_tail),
        .i_dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld(dp_lnk_cross_north_to_center_512_b_egr_rd_req_to_lnk_cross_north_to_center_512_b_ingr_rd_req_vld),
        .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_data),
        .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_head),
        .i_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld(dp_lnk_cross_north_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_north_to_center_512_b_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_data),
        .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_head),
        .o_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_rdy),
        .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_tail),
        .i_dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld(dp_lnk_cross_north_to_center_64_egr_req_to_lnk_cross_north_to_center_64_ingr_req_vld),
        .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_data),
        .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_head),
        .i_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_tail),
        .o_dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld(dp_lnk_cross_north_to_center_64_ingr_req_resp_to_lnk_cross_north_to_center_64_egr_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_data),
        .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_head),
        .o_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_tail),
        .i_dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_0_egr_rd_req_to_lnk_cross_south_to_center_512_0_ingr_rd_req_vld),
        .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_0_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_0_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_data),
        .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_head),
        .o_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_tail),
        .i_dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_1_egr_wr_req_to_lnk_cross_south_to_center_512_1_ingr_wr_req_vld),
        .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_1_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_1_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_data),
        .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_head),
        .o_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_tail),
        .i_dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_2_egr_wr_req_to_lnk_cross_south_to_center_512_2_ingr_wr_req_vld),
        .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_2_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_2_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_data),
        .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_head),
        .o_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_tail),
        .i_dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_3_egr_rd_req_to_lnk_cross_south_to_center_512_3_ingr_rd_req_vld),
        .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_3_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_3_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_data),
        .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_head),
        .o_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_tail),
        .i_dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_4_egr_rd_req_to_lnk_cross_south_to_center_512_4_ingr_rd_req_vld),
        .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_4_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_4_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_data),
        .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_head),
        .o_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_tail),
        .i_dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_5_egr_wr_req_to_lnk_cross_south_to_center_512_5_ingr_wr_req_vld),
        .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_5_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_5_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_data),
        .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_head),
        .o_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_tail),
        .i_dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_6_egr_wr_req_to_lnk_cross_south_to_center_512_6_ingr_wr_req_vld),
        .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_6_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_6_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_data),
        .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_head),
        .o_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_tail),
        .i_dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_7_egr_wr_req_to_lnk_cross_south_to_center_512_7_ingr_wr_req_vld),
        .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_7_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_7_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_data),
        .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_head),
        .o_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_tail),
        .i_dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_8_egr_rd_req_to_lnk_cross_south_to_center_512_8_ingr_rd_req_vld),
        .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_8_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_8_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_data),
        .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_head),
        .o_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_tail),
        .i_dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_9_egr_rd_req_to_lnk_cross_south_to_center_512_9_ingr_rd_req_vld),
        .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_9_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_9_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_data),
        .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_head),
        .o_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_tail),
        .i_dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld(dp_lnk_cross_south_to_center_512_a_egr_wr_req_to_lnk_cross_south_to_center_512_a_ingr_wr_req_vld),
        .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld(dp_lnk_cross_south_to_center_512_a_ingr_wr_req_resp_to_lnk_cross_south_to_center_512_a_egr_wr_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_data),
        .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_head),
        .o_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_rdy),
        .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_tail),
        .i_dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld(dp_lnk_cross_south_to_center_512_b_egr_rd_req_to_lnk_cross_south_to_center_512_b_ingr_rd_req_vld),
        .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_data),
        .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_head),
        .i_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld(dp_lnk_cross_south_to_center_512_b_ingr_rd_req_resp_to_lnk_cross_south_to_center_512_b_egr_rd_req_resp_vld),
        .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_data),
        .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_head),
        .o_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_rdy),
        .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_tail),
        .i_dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld(dp_lnk_cross_south_to_center_64_egr_req_to_lnk_cross_south_to_center_64_ingr_req_vld),
        .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_data),
        .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_head),
        .i_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_rdy),
        .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_tail),
        .o_dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld(dp_lnk_cross_south_to_center_64_ingr_req_resp_to_lnk_cross_south_to_center_64_egr_req_resp_vld),
        .i_l2_addr_mode_port_b0(i_l2_addr_mode_port_b0),
        .i_l2_addr_mode_port_b1(i_l2_addr_mode_port_b1),
        .i_l2_intr_mode_port_b0(i_l2_intr_mode_port_b0),
        .i_l2_intr_mode_port_b1(i_l2_intr_mode_port_b1),
        .i_lpddr_graph_addr_mode_port_b0(i_lpddr_graph_addr_mode_port_b0),
        .i_lpddr_graph_addr_mode_port_b1(i_lpddr_graph_addr_mode_port_b1),
        .i_lpddr_graph_intr_mode_port_b0(i_lpddr_graph_intr_mode_port_b0),
        .i_lpddr_graph_intr_mode_port_b1(i_lpddr_graph_intr_mode_port_b1),
        .i_lpddr_ppp_addr_mode_port_b0(i_lpddr_ppp_addr_mode_port_b0),
        .i_lpddr_ppp_addr_mode_port_b1(i_lpddr_ppp_addr_mode_port_b1),
        .i_lpddr_ppp_intr_mode_port_b0(i_lpddr_ppp_intr_mode_port_b0),
        .i_lpddr_ppp_intr_mode_port_b1(i_lpddr_ppp_intr_mode_port_b1),

        // Token Network IOs
        // - Fences
        .i_sdma_0_pwr_tok_idle_req(center_to_sdma_0_noc_tok_async_idle_req),
        .o_sdma_0_pwr_tok_idle_ack(center_to_sdma_0_noc_tok_async_idle_ack),
        .o_sdma_0_pwr_tok_idle_val(center_to_sdma_0_noc_tok_async_idle_val),
        .i_sdma_1_pwr_tok_idle_req(center_to_sdma_1_noc_tok_async_idle_req),
        .o_sdma_1_pwr_tok_idle_ack(center_to_sdma_1_noc_tok_async_idle_ack),
        .o_sdma_1_pwr_tok_idle_val(center_to_sdma_1_noc_tok_async_idle_val),

        // - NIUs
        .i_sdma_0_init_tok_ocpl_s_maddr     (sdma_0_init_tok_ocpl_maddr),
        .i_sdma_0_init_tok_ocpl_s_mcmd      (sdma_0_init_tok_ocpl_mcmd),
        .o_sdma_0_init_tok_ocpl_s_scmdaccept(sdma_0_init_tok_ocpl_scmdaccept),
        .i_sdma_0_init_tok_ocpl_s_mdata     (sdma_0_init_tok_ocpl_mdata),
        .o_sdma_0_targ_tok_ocpl_m_maddr     (sdma_0_targ_tok_ocpl_maddr),
        .o_sdma_0_targ_tok_ocpl_m_mcmd      (sdma_0_targ_tok_ocpl_mcmd),
        .i_sdma_0_targ_tok_ocpl_m_scmdaccept(sdma_0_targ_tok_ocpl_scmdaccept),
        .o_sdma_0_targ_tok_ocpl_m_mdata     (sdma_0_targ_tok_ocpl_mdata),
        .i_sdma_1_init_tok_ocpl_s_maddr     (sdma_1_init_tok_ocpl_maddr),
        .i_sdma_1_init_tok_ocpl_s_mcmd      (sdma_1_init_tok_ocpl_mcmd),
        .o_sdma_1_init_tok_ocpl_s_scmdaccept(sdma_1_init_tok_ocpl_scmdaccept),
        .i_sdma_1_init_tok_ocpl_s_mdata     (sdma_1_init_tok_ocpl_mdata),
        .o_sdma_1_targ_tok_ocpl_m_maddr     (sdma_1_targ_tok_ocpl_maddr),
        .o_sdma_1_targ_tok_ocpl_m_mcmd      (sdma_1_targ_tok_ocpl_mcmd),
        .i_sdma_1_targ_tok_ocpl_m_scmdaccept(sdma_1_targ_tok_ocpl_scmdaccept),
        .o_sdma_1_targ_tok_ocpl_m_mdata     (sdma_1_targ_tok_ocpl_mdata),

        .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_data),
        .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_head),
        .i_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_rdy),
        .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_tail),
        .o_dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld(dp_lnk_cross_center_to_east_tok_0_egress_to_lnk_cross_center_to_east_tok_0_ingress_vld),
        .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_data),
        .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_head),
        .i_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_rdy),
        .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_tail),
        .o_dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld(dp_lnk_cross_center_to_east_tok_1_egress_to_lnk_cross_center_to_east_tok_1_ingress_vld),
        .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_data),
        .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_head),
        .i_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_rdy),
        .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_tail),
        .o_dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld(dp_lnk_cross_center_to_north_tok_0_egress_to_lnk_cross_center_to_north_tok_0_ingress_vld),
        .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_data),
        .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_head),
        .i_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_rdy),
        .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_tail),
        .o_dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld(dp_lnk_cross_center_to_north_tok_1_egress_to_lnk_cross_center_to_north_tok_1_ingress_vld),
        .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_data),
        .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_head),
        .i_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_rdy),
        .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_tail),
        .o_dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld(dp_lnk_cross_center_to_south_tok_0_egress_to_lnk_cross_center_to_south_tok_0_ingress_vld),
        .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_data),
        .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_head),
        .i_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_rdy),
        .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_tail),
        .o_dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld(dp_lnk_cross_center_to_south_tok_1_egress_to_lnk_cross_center_to_south_tok_1_ingress_vld),
        .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_data),
        .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_head),
        .o_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_rdy),
        .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_tail),
        .i_dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld(dp_lnk_cross_east_to_center_tok_0_egress_to_lnk_cross_east_to_center_tok_0_ingress_vld),
        .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_data),
        .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_head),
        .o_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_rdy),
        .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_tail),
        .i_dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld(dp_lnk_cross_east_to_center_tok_1_egress_to_lnk_cross_east_to_center_tok_1_ingress_vld),
        .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_data),
        .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_head),
        .o_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_rdy),
        .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_tail),
        .i_dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld(dp_lnk_cross_north_to_center_tok_0_egress_to_lnk_cross_north_to_center_tok_0_ingress_vld),
        .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_data),
        .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_head),
        .o_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_rdy),
        .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_tail),
        .i_dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld(dp_lnk_cross_north_to_center_tok_1_egress_to_lnk_cross_north_to_center_tok_1_ingress_vld),
        .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_data),
        .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_head),
        .o_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_rdy),
        .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_tail),
        .i_dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld(dp_lnk_cross_south_to_center_tok_0_egress_to_lnk_cross_south_to_center_tok_0_ingress_vld),
        .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_data),
        .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_head),
        .o_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_rdy),
        .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_tail),
        .i_dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld(dp_lnk_cross_south_to_center_tok_1_egress_to_lnk_cross_south_to_center_tok_1_ingress_vld),

        .i_noc_clk(i_noc_clk),
        .i_noc_rst_n(i_noc_rst_n),
        .tck('0),
        .trst('0),
        .tms('0),
        .tdi('0),
        .tdo_en( ),
        .tdo( ),
        .test_clk('0),
        .test_mode(test_mode),
        .edt_update('0),
        .scan_en(scan_en),
        .scan_in('0),
        .scan_out(  )
    );
endmodule
