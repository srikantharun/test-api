
package lpddr_env_pkg;
  import lpddr_regs_pkg_uvm::*;
  
  `include "subsystem_signal_intf.sv"

endpackage : lpddr_env_pkg
